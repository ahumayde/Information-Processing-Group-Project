// esp32SPIHardware.v

// Generated using ACDS version 20.1 711

`timescale 1 ps / 1 ps
module esp32SPIHardware (
		inout  wire        accelerometer_spi_I2C_SDAT,      // accelerometer_spi.I2C_SDAT
		output wire        accelerometer_spi_I2C_SCLK,      //                  .I2C_SCLK
		output wire        accelerometer_spi_G_SENSOR_CS_N, //                  .G_SENSOR_CS_N
		input  wire        accelerometer_spi_G_SENSOR_INT,  //                  .G_SENSOR_INT
		input  wire        clk_clk,                         //               clk.clk
		output wire [12:0] dram_addr,                       //              dram.addr
		output wire [1:0]  dram_ba,                         //                  .ba
		output wire        dram_cas_n,                      //                  .cas_n
		output wire        dram_cke,                        //                  .cke
		output wire        dram_cs_n,                       //                  .cs_n
		inout  wire [15:0] dram_dq,                         //                  .dq
		output wire [1:0]  dram_dqm,                        //                  .dqm
		output wire        dram_ras_n,                      //                  .ras_n
		output wire        dram_we_n,                       //                  .we_n
		input  wire        esp32_spi_MISO,                  //         esp32_spi.MISO
		output wire        esp32_spi_MOSI,                  //                  .MOSI
		output wire        esp32_spi_SCLK,                  //                  .SCLK
		output wire        esp32_spi_SS_n,                  //                  .SS_n
		input  wire        reset_reset_n,                   //             reset.reset_n
		output wire        sdram_clk_clk                    //         sdram_clk.clk
	);

	wire         dram_clks_pll_sys_clk_clk;                                                       // dram_clks_pll:sys_clk_clk -> [accelerometer:clk, dram_controller:clk, esp32_spi:clk, irq_mapper:clk, jtag:clk, mm_interconnect_0:dram_clks_pll_sys_clk_clk, nios2_cpu:clk, rst_controller:clk, sys_clk:clk, timer_1:clk, timer_2:clk]
	wire         nios2_cpu_custom_instruction_master_readra;                                      // nios2_cpu:E_ci_combo_readra -> nios2_cpu_custom_instruction_master_translator:ci_slave_readra
	wire         nios2_cpu_custom_instruction_master_readrb;                                      // nios2_cpu:E_ci_combo_readrb -> nios2_cpu_custom_instruction_master_translator:ci_slave_readrb
	wire   [4:0] nios2_cpu_custom_instruction_master_multi_b;                                     // nios2_cpu:A_ci_multi_b -> nios2_cpu_custom_instruction_master_translator:ci_slave_multi_b
	wire   [4:0] nios2_cpu_custom_instruction_master_multi_c;                                     // nios2_cpu:A_ci_multi_c -> nios2_cpu_custom_instruction_master_translator:ci_slave_multi_c
	wire         nios2_cpu_custom_instruction_master_reset_req;                                   // nios2_cpu:A_ci_multi_reset_req -> nios2_cpu_custom_instruction_master_translator:ci_slave_multi_reset_req
	wire   [4:0] nios2_cpu_custom_instruction_master_multi_a;                                     // nios2_cpu:A_ci_multi_a -> nios2_cpu_custom_instruction_master_translator:ci_slave_multi_a
	wire  [31:0] nios2_cpu_custom_instruction_master_result;                                      // nios2_cpu_custom_instruction_master_translator:ci_slave_result -> nios2_cpu:E_ci_combo_result
	wire  [31:0] nios2_cpu_custom_instruction_master_datab;                                       // nios2_cpu:E_ci_combo_datab -> nios2_cpu_custom_instruction_master_translator:ci_slave_datab
	wire  [31:0] nios2_cpu_custom_instruction_master_dataa;                                       // nios2_cpu:E_ci_combo_dataa -> nios2_cpu_custom_instruction_master_translator:ci_slave_dataa
	wire         nios2_cpu_custom_instruction_master_writerc;                                     // nios2_cpu:E_ci_combo_writerc -> nios2_cpu_custom_instruction_master_translator:ci_slave_writerc
	wire  [31:0] nios2_cpu_custom_instruction_master_multi_dataa;                                 // nios2_cpu:A_ci_multi_dataa -> nios2_cpu_custom_instruction_master_translator:ci_slave_multi_dataa
	wire         nios2_cpu_custom_instruction_master_multi_writerc;                               // nios2_cpu:A_ci_multi_writerc -> nios2_cpu_custom_instruction_master_translator:ci_slave_multi_writerc
	wire   [4:0] nios2_cpu_custom_instruction_master_a;                                           // nios2_cpu:E_ci_combo_a -> nios2_cpu_custom_instruction_master_translator:ci_slave_a
	wire   [4:0] nios2_cpu_custom_instruction_master_b;                                           // nios2_cpu:E_ci_combo_b -> nios2_cpu_custom_instruction_master_translator:ci_slave_b
	wire  [31:0] nios2_cpu_custom_instruction_master_multi_result;                                // nios2_cpu_custom_instruction_master_translator:ci_slave_multi_result -> nios2_cpu:A_ci_multi_result
	wire         nios2_cpu_custom_instruction_master_clk;                                         // nios2_cpu:A_ci_multi_clock -> nios2_cpu_custom_instruction_master_translator:ci_slave_multi_clk
	wire  [31:0] nios2_cpu_custom_instruction_master_multi_datab;                                 // nios2_cpu:A_ci_multi_datab -> nios2_cpu_custom_instruction_master_translator:ci_slave_multi_datab
	wire   [4:0] nios2_cpu_custom_instruction_master_c;                                           // nios2_cpu:E_ci_combo_c -> nios2_cpu_custom_instruction_master_translator:ci_slave_c
	wire  [31:0] nios2_cpu_custom_instruction_master_ipending;                                    // nios2_cpu:E_ci_combo_ipending -> nios2_cpu_custom_instruction_master_translator:ci_slave_ipending
	wire         nios2_cpu_custom_instruction_master_start;                                       // nios2_cpu:A_ci_multi_start -> nios2_cpu_custom_instruction_master_translator:ci_slave_multi_start
	wire         nios2_cpu_custom_instruction_master_done;                                        // nios2_cpu_custom_instruction_master_translator:ci_slave_multi_done -> nios2_cpu:A_ci_multi_done
	wire   [7:0] nios2_cpu_custom_instruction_master_n;                                           // nios2_cpu:E_ci_combo_n -> nios2_cpu_custom_instruction_master_translator:ci_slave_n
	wire         nios2_cpu_custom_instruction_master_estatus;                                     // nios2_cpu:E_ci_combo_estatus -> nios2_cpu_custom_instruction_master_translator:ci_slave_estatus
	wire         nios2_cpu_custom_instruction_master_clk_en;                                      // nios2_cpu:A_ci_multi_clk_en -> nios2_cpu_custom_instruction_master_translator:ci_slave_multi_clken
	wire         nios2_cpu_custom_instruction_master_reset;                                       // nios2_cpu:A_ci_multi_reset -> nios2_cpu_custom_instruction_master_translator:ci_slave_multi_reset
	wire         nios2_cpu_custom_instruction_master_multi_readrb;                                // nios2_cpu:A_ci_multi_readrb -> nios2_cpu_custom_instruction_master_translator:ci_slave_multi_readrb
	wire         nios2_cpu_custom_instruction_master_multi_readra;                                // nios2_cpu:A_ci_multi_readra -> nios2_cpu_custom_instruction_master_translator:ci_slave_multi_readra
	wire   [7:0] nios2_cpu_custom_instruction_master_multi_n;                                     // nios2_cpu:A_ci_multi_n -> nios2_cpu_custom_instruction_master_translator:ci_slave_multi_n
	wire  [31:0] nios2_cpu_custom_instruction_master_translator_comb_ci_master_result;            // nios2_cpu_custom_instruction_master_comb_xconnect:ci_slave_result -> nios2_cpu_custom_instruction_master_translator:comb_ci_master_result
	wire         nios2_cpu_custom_instruction_master_translator_comb_ci_master_readra;            // nios2_cpu_custom_instruction_master_translator:comb_ci_master_readra -> nios2_cpu_custom_instruction_master_comb_xconnect:ci_slave_readra
	wire   [4:0] nios2_cpu_custom_instruction_master_translator_comb_ci_master_a;                 // nios2_cpu_custom_instruction_master_translator:comb_ci_master_a -> nios2_cpu_custom_instruction_master_comb_xconnect:ci_slave_a
	wire   [4:0] nios2_cpu_custom_instruction_master_translator_comb_ci_master_b;                 // nios2_cpu_custom_instruction_master_translator:comb_ci_master_b -> nios2_cpu_custom_instruction_master_comb_xconnect:ci_slave_b
	wire         nios2_cpu_custom_instruction_master_translator_comb_ci_master_readrb;            // nios2_cpu_custom_instruction_master_translator:comb_ci_master_readrb -> nios2_cpu_custom_instruction_master_comb_xconnect:ci_slave_readrb
	wire   [4:0] nios2_cpu_custom_instruction_master_translator_comb_ci_master_c;                 // nios2_cpu_custom_instruction_master_translator:comb_ci_master_c -> nios2_cpu_custom_instruction_master_comb_xconnect:ci_slave_c
	wire         nios2_cpu_custom_instruction_master_translator_comb_ci_master_estatus;           // nios2_cpu_custom_instruction_master_translator:comb_ci_master_estatus -> nios2_cpu_custom_instruction_master_comb_xconnect:ci_slave_estatus
	wire  [31:0] nios2_cpu_custom_instruction_master_translator_comb_ci_master_ipending;          // nios2_cpu_custom_instruction_master_translator:comb_ci_master_ipending -> nios2_cpu_custom_instruction_master_comb_xconnect:ci_slave_ipending
	wire  [31:0] nios2_cpu_custom_instruction_master_translator_comb_ci_master_datab;             // nios2_cpu_custom_instruction_master_translator:comb_ci_master_datab -> nios2_cpu_custom_instruction_master_comb_xconnect:ci_slave_datab
	wire  [31:0] nios2_cpu_custom_instruction_master_translator_comb_ci_master_dataa;             // nios2_cpu_custom_instruction_master_translator:comb_ci_master_dataa -> nios2_cpu_custom_instruction_master_comb_xconnect:ci_slave_dataa
	wire         nios2_cpu_custom_instruction_master_translator_comb_ci_master_writerc;           // nios2_cpu_custom_instruction_master_translator:comb_ci_master_writerc -> nios2_cpu_custom_instruction_master_comb_xconnect:ci_slave_writerc
	wire   [7:0] nios2_cpu_custom_instruction_master_translator_comb_ci_master_n;                 // nios2_cpu_custom_instruction_master_translator:comb_ci_master_n -> nios2_cpu_custom_instruction_master_comb_xconnect:ci_slave_n
	wire  [31:0] nios2_cpu_custom_instruction_master_comb_xconnect_ci_master0_result;             // nios2_cpu_custom_instruction_master_comb_slave_translator0:ci_slave_result -> nios2_cpu_custom_instruction_master_comb_xconnect:ci_master0_result
	wire         nios2_cpu_custom_instruction_master_comb_xconnect_ci_master0_readra;             // nios2_cpu_custom_instruction_master_comb_xconnect:ci_master0_readra -> nios2_cpu_custom_instruction_master_comb_slave_translator0:ci_slave_readra
	wire   [4:0] nios2_cpu_custom_instruction_master_comb_xconnect_ci_master0_a;                  // nios2_cpu_custom_instruction_master_comb_xconnect:ci_master0_a -> nios2_cpu_custom_instruction_master_comb_slave_translator0:ci_slave_a
	wire   [4:0] nios2_cpu_custom_instruction_master_comb_xconnect_ci_master0_b;                  // nios2_cpu_custom_instruction_master_comb_xconnect:ci_master0_b -> nios2_cpu_custom_instruction_master_comb_slave_translator0:ci_slave_b
	wire         nios2_cpu_custom_instruction_master_comb_xconnect_ci_master0_readrb;             // nios2_cpu_custom_instruction_master_comb_xconnect:ci_master0_readrb -> nios2_cpu_custom_instruction_master_comb_slave_translator0:ci_slave_readrb
	wire   [4:0] nios2_cpu_custom_instruction_master_comb_xconnect_ci_master0_c;                  // nios2_cpu_custom_instruction_master_comb_xconnect:ci_master0_c -> nios2_cpu_custom_instruction_master_comb_slave_translator0:ci_slave_c
	wire         nios2_cpu_custom_instruction_master_comb_xconnect_ci_master0_estatus;            // nios2_cpu_custom_instruction_master_comb_xconnect:ci_master0_estatus -> nios2_cpu_custom_instruction_master_comb_slave_translator0:ci_slave_estatus
	wire  [31:0] nios2_cpu_custom_instruction_master_comb_xconnect_ci_master0_ipending;           // nios2_cpu_custom_instruction_master_comb_xconnect:ci_master0_ipending -> nios2_cpu_custom_instruction_master_comb_slave_translator0:ci_slave_ipending
	wire  [31:0] nios2_cpu_custom_instruction_master_comb_xconnect_ci_master0_datab;              // nios2_cpu_custom_instruction_master_comb_xconnect:ci_master0_datab -> nios2_cpu_custom_instruction_master_comb_slave_translator0:ci_slave_datab
	wire  [31:0] nios2_cpu_custom_instruction_master_comb_xconnect_ci_master0_dataa;              // nios2_cpu_custom_instruction_master_comb_xconnect:ci_master0_dataa -> nios2_cpu_custom_instruction_master_comb_slave_translator0:ci_slave_dataa
	wire         nios2_cpu_custom_instruction_master_comb_xconnect_ci_master0_writerc;            // nios2_cpu_custom_instruction_master_comb_xconnect:ci_master0_writerc -> nios2_cpu_custom_instruction_master_comb_slave_translator0:ci_slave_writerc
	wire   [7:0] nios2_cpu_custom_instruction_master_comb_xconnect_ci_master0_n;                  // nios2_cpu_custom_instruction_master_comb_xconnect:ci_master0_n -> nios2_cpu_custom_instruction_master_comb_slave_translator0:ci_slave_n
	wire  [31:0] nios2_cpu_custom_instruction_master_comb_slave_translator0_ci_master_result;     // fph2:s1_result -> nios2_cpu_custom_instruction_master_comb_slave_translator0:ci_master_result
	wire  [31:0] nios2_cpu_custom_instruction_master_comb_slave_translator0_ci_master_datab;      // nios2_cpu_custom_instruction_master_comb_slave_translator0:ci_master_datab -> fph2:s1_datab
	wire  [31:0] nios2_cpu_custom_instruction_master_comb_slave_translator0_ci_master_dataa;      // nios2_cpu_custom_instruction_master_comb_slave_translator0:ci_master_dataa -> fph2:s1_dataa
	wire   [3:0] nios2_cpu_custom_instruction_master_comb_slave_translator0_ci_master_n;          // nios2_cpu_custom_instruction_master_comb_slave_translator0:ci_master_n -> fph2:s1_n
	wire         nios2_cpu_custom_instruction_master_translator_multi_ci_master_readra;           // nios2_cpu_custom_instruction_master_translator:multi_ci_master_readra -> nios2_cpu_custom_instruction_master_multi_xconnect:ci_slave_readra
	wire   [4:0] nios2_cpu_custom_instruction_master_translator_multi_ci_master_a;                // nios2_cpu_custom_instruction_master_translator:multi_ci_master_a -> nios2_cpu_custom_instruction_master_multi_xconnect:ci_slave_a
	wire   [4:0] nios2_cpu_custom_instruction_master_translator_multi_ci_master_b;                // nios2_cpu_custom_instruction_master_translator:multi_ci_master_b -> nios2_cpu_custom_instruction_master_multi_xconnect:ci_slave_b
	wire         nios2_cpu_custom_instruction_master_translator_multi_ci_master_clk;              // nios2_cpu_custom_instruction_master_translator:multi_ci_master_clk -> nios2_cpu_custom_instruction_master_multi_xconnect:ci_slave_clk
	wire         nios2_cpu_custom_instruction_master_translator_multi_ci_master_readrb;           // nios2_cpu_custom_instruction_master_translator:multi_ci_master_readrb -> nios2_cpu_custom_instruction_master_multi_xconnect:ci_slave_readrb
	wire   [4:0] nios2_cpu_custom_instruction_master_translator_multi_ci_master_c;                // nios2_cpu_custom_instruction_master_translator:multi_ci_master_c -> nios2_cpu_custom_instruction_master_multi_xconnect:ci_slave_c
	wire         nios2_cpu_custom_instruction_master_translator_multi_ci_master_start;            // nios2_cpu_custom_instruction_master_translator:multi_ci_master_start -> nios2_cpu_custom_instruction_master_multi_xconnect:ci_slave_start
	wire         nios2_cpu_custom_instruction_master_translator_multi_ci_master_reset_req;        // nios2_cpu_custom_instruction_master_translator:multi_ci_master_reset_req -> nios2_cpu_custom_instruction_master_multi_xconnect:ci_slave_reset_req
	wire         nios2_cpu_custom_instruction_master_translator_multi_ci_master_done;             // nios2_cpu_custom_instruction_master_multi_xconnect:ci_slave_done -> nios2_cpu_custom_instruction_master_translator:multi_ci_master_done
	wire   [7:0] nios2_cpu_custom_instruction_master_translator_multi_ci_master_n;                // nios2_cpu_custom_instruction_master_translator:multi_ci_master_n -> nios2_cpu_custom_instruction_master_multi_xconnect:ci_slave_n
	wire  [31:0] nios2_cpu_custom_instruction_master_translator_multi_ci_master_result;           // nios2_cpu_custom_instruction_master_multi_xconnect:ci_slave_result -> nios2_cpu_custom_instruction_master_translator:multi_ci_master_result
	wire         nios2_cpu_custom_instruction_master_translator_multi_ci_master_clk_en;           // nios2_cpu_custom_instruction_master_translator:multi_ci_master_clken -> nios2_cpu_custom_instruction_master_multi_xconnect:ci_slave_clken
	wire  [31:0] nios2_cpu_custom_instruction_master_translator_multi_ci_master_datab;            // nios2_cpu_custom_instruction_master_translator:multi_ci_master_datab -> nios2_cpu_custom_instruction_master_multi_xconnect:ci_slave_datab
	wire  [31:0] nios2_cpu_custom_instruction_master_translator_multi_ci_master_dataa;            // nios2_cpu_custom_instruction_master_translator:multi_ci_master_dataa -> nios2_cpu_custom_instruction_master_multi_xconnect:ci_slave_dataa
	wire         nios2_cpu_custom_instruction_master_translator_multi_ci_master_reset;            // nios2_cpu_custom_instruction_master_translator:multi_ci_master_reset -> nios2_cpu_custom_instruction_master_multi_xconnect:ci_slave_reset
	wire         nios2_cpu_custom_instruction_master_translator_multi_ci_master_writerc;          // nios2_cpu_custom_instruction_master_translator:multi_ci_master_writerc -> nios2_cpu_custom_instruction_master_multi_xconnect:ci_slave_writerc
	wire         nios2_cpu_custom_instruction_master_multi_xconnect_ci_master0_readra;            // nios2_cpu_custom_instruction_master_multi_xconnect:ci_master0_readra -> nios2_cpu_custom_instruction_master_multi_slave_translator0:ci_slave_readra
	wire   [4:0] nios2_cpu_custom_instruction_master_multi_xconnect_ci_master0_a;                 // nios2_cpu_custom_instruction_master_multi_xconnect:ci_master0_a -> nios2_cpu_custom_instruction_master_multi_slave_translator0:ci_slave_a
	wire   [4:0] nios2_cpu_custom_instruction_master_multi_xconnect_ci_master0_b;                 // nios2_cpu_custom_instruction_master_multi_xconnect:ci_master0_b -> nios2_cpu_custom_instruction_master_multi_slave_translator0:ci_slave_b
	wire         nios2_cpu_custom_instruction_master_multi_xconnect_ci_master0_readrb;            // nios2_cpu_custom_instruction_master_multi_xconnect:ci_master0_readrb -> nios2_cpu_custom_instruction_master_multi_slave_translator0:ci_slave_readrb
	wire   [4:0] nios2_cpu_custom_instruction_master_multi_xconnect_ci_master0_c;                 // nios2_cpu_custom_instruction_master_multi_xconnect:ci_master0_c -> nios2_cpu_custom_instruction_master_multi_slave_translator0:ci_slave_c
	wire         nios2_cpu_custom_instruction_master_multi_xconnect_ci_master0_clk;               // nios2_cpu_custom_instruction_master_multi_xconnect:ci_master0_clk -> nios2_cpu_custom_instruction_master_multi_slave_translator0:ci_slave_clk
	wire  [31:0] nios2_cpu_custom_instruction_master_multi_xconnect_ci_master0_ipending;          // nios2_cpu_custom_instruction_master_multi_xconnect:ci_master0_ipending -> nios2_cpu_custom_instruction_master_multi_slave_translator0:ci_slave_ipending
	wire         nios2_cpu_custom_instruction_master_multi_xconnect_ci_master0_start;             // nios2_cpu_custom_instruction_master_multi_xconnect:ci_master0_start -> nios2_cpu_custom_instruction_master_multi_slave_translator0:ci_slave_start
	wire         nios2_cpu_custom_instruction_master_multi_xconnect_ci_master0_reset_req;         // nios2_cpu_custom_instruction_master_multi_xconnect:ci_master0_reset_req -> nios2_cpu_custom_instruction_master_multi_slave_translator0:ci_slave_reset_req
	wire         nios2_cpu_custom_instruction_master_multi_xconnect_ci_master0_done;              // nios2_cpu_custom_instruction_master_multi_slave_translator0:ci_slave_done -> nios2_cpu_custom_instruction_master_multi_xconnect:ci_master0_done
	wire   [7:0] nios2_cpu_custom_instruction_master_multi_xconnect_ci_master0_n;                 // nios2_cpu_custom_instruction_master_multi_xconnect:ci_master0_n -> nios2_cpu_custom_instruction_master_multi_slave_translator0:ci_slave_n
	wire  [31:0] nios2_cpu_custom_instruction_master_multi_xconnect_ci_master0_result;            // nios2_cpu_custom_instruction_master_multi_slave_translator0:ci_slave_result -> nios2_cpu_custom_instruction_master_multi_xconnect:ci_master0_result
	wire         nios2_cpu_custom_instruction_master_multi_xconnect_ci_master0_estatus;           // nios2_cpu_custom_instruction_master_multi_xconnect:ci_master0_estatus -> nios2_cpu_custom_instruction_master_multi_slave_translator0:ci_slave_estatus
	wire         nios2_cpu_custom_instruction_master_multi_xconnect_ci_master0_clk_en;            // nios2_cpu_custom_instruction_master_multi_xconnect:ci_master0_clken -> nios2_cpu_custom_instruction_master_multi_slave_translator0:ci_slave_clken
	wire  [31:0] nios2_cpu_custom_instruction_master_multi_xconnect_ci_master0_datab;             // nios2_cpu_custom_instruction_master_multi_xconnect:ci_master0_datab -> nios2_cpu_custom_instruction_master_multi_slave_translator0:ci_slave_datab
	wire  [31:0] nios2_cpu_custom_instruction_master_multi_xconnect_ci_master0_dataa;             // nios2_cpu_custom_instruction_master_multi_xconnect:ci_master0_dataa -> nios2_cpu_custom_instruction_master_multi_slave_translator0:ci_slave_dataa
	wire         nios2_cpu_custom_instruction_master_multi_xconnect_ci_master0_reset;             // nios2_cpu_custom_instruction_master_multi_xconnect:ci_master0_reset -> nios2_cpu_custom_instruction_master_multi_slave_translator0:ci_slave_reset
	wire         nios2_cpu_custom_instruction_master_multi_xconnect_ci_master0_writerc;           // nios2_cpu_custom_instruction_master_multi_xconnect:ci_master0_writerc -> nios2_cpu_custom_instruction_master_multi_slave_translator0:ci_slave_writerc
	wire  [31:0] nios2_cpu_custom_instruction_master_multi_slave_translator0_ci_master_result;    // fph2:s2_result -> nios2_cpu_custom_instruction_master_multi_slave_translator0:ci_master_result
	wire         nios2_cpu_custom_instruction_master_multi_slave_translator0_ci_master_clk;       // nios2_cpu_custom_instruction_master_multi_slave_translator0:ci_master_clk -> fph2:s2_clk
	wire         nios2_cpu_custom_instruction_master_multi_slave_translator0_ci_master_clk_en;    // nios2_cpu_custom_instruction_master_multi_slave_translator0:ci_master_clken -> fph2:s2_clk_en
	wire  [31:0] nios2_cpu_custom_instruction_master_multi_slave_translator0_ci_master_datab;     // nios2_cpu_custom_instruction_master_multi_slave_translator0:ci_master_datab -> fph2:s2_datab
	wire  [31:0] nios2_cpu_custom_instruction_master_multi_slave_translator0_ci_master_dataa;     // nios2_cpu_custom_instruction_master_multi_slave_translator0:ci_master_dataa -> fph2:s2_dataa
	wire         nios2_cpu_custom_instruction_master_multi_slave_translator0_ci_master_start;     // nios2_cpu_custom_instruction_master_multi_slave_translator0:ci_master_start -> fph2:s2_start
	wire         nios2_cpu_custom_instruction_master_multi_slave_translator0_ci_master_reset;     // nios2_cpu_custom_instruction_master_multi_slave_translator0:ci_master_reset -> fph2:s2_reset
	wire         nios2_cpu_custom_instruction_master_multi_slave_translator0_ci_master_reset_req; // nios2_cpu_custom_instruction_master_multi_slave_translator0:ci_master_reset_req -> fph2:s2_reset_req
	wire         nios2_cpu_custom_instruction_master_multi_slave_translator0_ci_master_done;      // fph2:s2_done -> nios2_cpu_custom_instruction_master_multi_slave_translator0:ci_master_done
	wire   [2:0] nios2_cpu_custom_instruction_master_multi_slave_translator0_ci_master_n;         // nios2_cpu_custom_instruction_master_multi_slave_translator0:ci_master_n -> fph2:s2_n
	wire  [31:0] nios2_cpu_data_master_readdata;                                                  // mm_interconnect_0:nios2_cpu_data_master_readdata -> nios2_cpu:d_readdata
	wire         nios2_cpu_data_master_waitrequest;                                               // mm_interconnect_0:nios2_cpu_data_master_waitrequest -> nios2_cpu:d_waitrequest
	wire         nios2_cpu_data_master_debugaccess;                                               // nios2_cpu:debug_mem_slave_debugaccess_to_roms -> mm_interconnect_0:nios2_cpu_data_master_debugaccess
	wire  [27:0] nios2_cpu_data_master_address;                                                   // nios2_cpu:d_address -> mm_interconnect_0:nios2_cpu_data_master_address
	wire   [3:0] nios2_cpu_data_master_byteenable;                                                // nios2_cpu:d_byteenable -> mm_interconnect_0:nios2_cpu_data_master_byteenable
	wire         nios2_cpu_data_master_read;                                                      // nios2_cpu:d_read -> mm_interconnect_0:nios2_cpu_data_master_read
	wire         nios2_cpu_data_master_readdatavalid;                                             // mm_interconnect_0:nios2_cpu_data_master_readdatavalid -> nios2_cpu:d_readdatavalid
	wire         nios2_cpu_data_master_write;                                                     // nios2_cpu:d_write -> mm_interconnect_0:nios2_cpu_data_master_write
	wire  [31:0] nios2_cpu_data_master_writedata;                                                 // nios2_cpu:d_writedata -> mm_interconnect_0:nios2_cpu_data_master_writedata
	wire  [31:0] nios2_cpu_instruction_master_readdata;                                           // mm_interconnect_0:nios2_cpu_instruction_master_readdata -> nios2_cpu:i_readdata
	wire         nios2_cpu_instruction_master_waitrequest;                                        // mm_interconnect_0:nios2_cpu_instruction_master_waitrequest -> nios2_cpu:i_waitrequest
	wire  [27:0] nios2_cpu_instruction_master_address;                                            // nios2_cpu:i_address -> mm_interconnect_0:nios2_cpu_instruction_master_address
	wire         nios2_cpu_instruction_master_read;                                               // nios2_cpu:i_read -> mm_interconnect_0:nios2_cpu_instruction_master_read
	wire         nios2_cpu_instruction_master_readdatavalid;                                      // mm_interconnect_0:nios2_cpu_instruction_master_readdatavalid -> nios2_cpu:i_readdatavalid
	wire   [7:0] mm_interconnect_0_accelerometer_avalon_accelerometer_spi_mode_slave_readdata;    // accelerometer:readdata -> mm_interconnect_0:accelerometer_avalon_accelerometer_spi_mode_slave_readdata
	wire         mm_interconnect_0_accelerometer_avalon_accelerometer_spi_mode_slave_waitrequest; // accelerometer:waitrequest -> mm_interconnect_0:accelerometer_avalon_accelerometer_spi_mode_slave_waitrequest
	wire   [0:0] mm_interconnect_0_accelerometer_avalon_accelerometer_spi_mode_slave_address;     // mm_interconnect_0:accelerometer_avalon_accelerometer_spi_mode_slave_address -> accelerometer:address
	wire         mm_interconnect_0_accelerometer_avalon_accelerometer_spi_mode_slave_read;        // mm_interconnect_0:accelerometer_avalon_accelerometer_spi_mode_slave_read -> accelerometer:read
	wire   [0:0] mm_interconnect_0_accelerometer_avalon_accelerometer_spi_mode_slave_byteenable;  // mm_interconnect_0:accelerometer_avalon_accelerometer_spi_mode_slave_byteenable -> accelerometer:byteenable
	wire         mm_interconnect_0_accelerometer_avalon_accelerometer_spi_mode_slave_write;       // mm_interconnect_0:accelerometer_avalon_accelerometer_spi_mode_slave_write -> accelerometer:write
	wire   [7:0] mm_interconnect_0_accelerometer_avalon_accelerometer_spi_mode_slave_writedata;   // mm_interconnect_0:accelerometer_avalon_accelerometer_spi_mode_slave_writedata -> accelerometer:writedata
	wire         mm_interconnect_0_jtag_avalon_jtag_slave_chipselect;                             // mm_interconnect_0:jtag_avalon_jtag_slave_chipselect -> jtag:av_chipselect
	wire  [31:0] mm_interconnect_0_jtag_avalon_jtag_slave_readdata;                               // jtag:av_readdata -> mm_interconnect_0:jtag_avalon_jtag_slave_readdata
	wire         mm_interconnect_0_jtag_avalon_jtag_slave_waitrequest;                            // jtag:av_waitrequest -> mm_interconnect_0:jtag_avalon_jtag_slave_waitrequest
	wire   [0:0] mm_interconnect_0_jtag_avalon_jtag_slave_address;                                // mm_interconnect_0:jtag_avalon_jtag_slave_address -> jtag:av_address
	wire         mm_interconnect_0_jtag_avalon_jtag_slave_read;                                   // mm_interconnect_0:jtag_avalon_jtag_slave_read -> jtag:av_read_n
	wire         mm_interconnect_0_jtag_avalon_jtag_slave_write;                                  // mm_interconnect_0:jtag_avalon_jtag_slave_write -> jtag:av_write_n
	wire  [31:0] mm_interconnect_0_jtag_avalon_jtag_slave_writedata;                              // mm_interconnect_0:jtag_avalon_jtag_slave_writedata -> jtag:av_writedata
	wire  [31:0] mm_interconnect_0_nios2_cpu_debug_mem_slave_readdata;                            // nios2_cpu:debug_mem_slave_readdata -> mm_interconnect_0:nios2_cpu_debug_mem_slave_readdata
	wire         mm_interconnect_0_nios2_cpu_debug_mem_slave_waitrequest;                         // nios2_cpu:debug_mem_slave_waitrequest -> mm_interconnect_0:nios2_cpu_debug_mem_slave_waitrequest
	wire         mm_interconnect_0_nios2_cpu_debug_mem_slave_debugaccess;                         // mm_interconnect_0:nios2_cpu_debug_mem_slave_debugaccess -> nios2_cpu:debug_mem_slave_debugaccess
	wire   [8:0] mm_interconnect_0_nios2_cpu_debug_mem_slave_address;                             // mm_interconnect_0:nios2_cpu_debug_mem_slave_address -> nios2_cpu:debug_mem_slave_address
	wire         mm_interconnect_0_nios2_cpu_debug_mem_slave_read;                                // mm_interconnect_0:nios2_cpu_debug_mem_slave_read -> nios2_cpu:debug_mem_slave_read
	wire   [3:0] mm_interconnect_0_nios2_cpu_debug_mem_slave_byteenable;                          // mm_interconnect_0:nios2_cpu_debug_mem_slave_byteenable -> nios2_cpu:debug_mem_slave_byteenable
	wire         mm_interconnect_0_nios2_cpu_debug_mem_slave_write;                               // mm_interconnect_0:nios2_cpu_debug_mem_slave_write -> nios2_cpu:debug_mem_slave_write
	wire  [31:0] mm_interconnect_0_nios2_cpu_debug_mem_slave_writedata;                           // mm_interconnect_0:nios2_cpu_debug_mem_slave_writedata -> nios2_cpu:debug_mem_slave_writedata
	wire         mm_interconnect_0_dram_controller_s1_chipselect;                                 // mm_interconnect_0:dram_controller_s1_chipselect -> dram_controller:az_cs
	wire  [15:0] mm_interconnect_0_dram_controller_s1_readdata;                                   // dram_controller:za_data -> mm_interconnect_0:dram_controller_s1_readdata
	wire         mm_interconnect_0_dram_controller_s1_waitrequest;                                // dram_controller:za_waitrequest -> mm_interconnect_0:dram_controller_s1_waitrequest
	wire  [24:0] mm_interconnect_0_dram_controller_s1_address;                                    // mm_interconnect_0:dram_controller_s1_address -> dram_controller:az_addr
	wire         mm_interconnect_0_dram_controller_s1_read;                                       // mm_interconnect_0:dram_controller_s1_read -> dram_controller:az_rd_n
	wire   [1:0] mm_interconnect_0_dram_controller_s1_byteenable;                                 // mm_interconnect_0:dram_controller_s1_byteenable -> dram_controller:az_be_n
	wire         mm_interconnect_0_dram_controller_s1_readdatavalid;                              // dram_controller:za_valid -> mm_interconnect_0:dram_controller_s1_readdatavalid
	wire         mm_interconnect_0_dram_controller_s1_write;                                      // mm_interconnect_0:dram_controller_s1_write -> dram_controller:az_wr_n
	wire  [15:0] mm_interconnect_0_dram_controller_s1_writedata;                                  // mm_interconnect_0:dram_controller_s1_writedata -> dram_controller:az_data
	wire         mm_interconnect_0_sys_clk_s1_chipselect;                                         // mm_interconnect_0:sys_clk_s1_chipselect -> sys_clk:chipselect
	wire  [15:0] mm_interconnect_0_sys_clk_s1_readdata;                                           // sys_clk:readdata -> mm_interconnect_0:sys_clk_s1_readdata
	wire   [2:0] mm_interconnect_0_sys_clk_s1_address;                                            // mm_interconnect_0:sys_clk_s1_address -> sys_clk:address
	wire         mm_interconnect_0_sys_clk_s1_write;                                              // mm_interconnect_0:sys_clk_s1_write -> sys_clk:write_n
	wire  [15:0] mm_interconnect_0_sys_clk_s1_writedata;                                          // mm_interconnect_0:sys_clk_s1_writedata -> sys_clk:writedata
	wire         mm_interconnect_0_timer_1_s1_chipselect;                                         // mm_interconnect_0:timer_1_s1_chipselect -> timer_1:chipselect
	wire  [15:0] mm_interconnect_0_timer_1_s1_readdata;                                           // timer_1:readdata -> mm_interconnect_0:timer_1_s1_readdata
	wire   [2:0] mm_interconnect_0_timer_1_s1_address;                                            // mm_interconnect_0:timer_1_s1_address -> timer_1:address
	wire         mm_interconnect_0_timer_1_s1_write;                                              // mm_interconnect_0:timer_1_s1_write -> timer_1:write_n
	wire  [15:0] mm_interconnect_0_timer_1_s1_writedata;                                          // mm_interconnect_0:timer_1_s1_writedata -> timer_1:writedata
	wire         mm_interconnect_0_timer_2_s1_chipselect;                                         // mm_interconnect_0:timer_2_s1_chipselect -> timer_2:chipselect
	wire  [15:0] mm_interconnect_0_timer_2_s1_readdata;                                           // timer_2:readdata -> mm_interconnect_0:timer_2_s1_readdata
	wire   [2:0] mm_interconnect_0_timer_2_s1_address;                                            // mm_interconnect_0:timer_2_s1_address -> timer_2:address
	wire         mm_interconnect_0_timer_2_s1_write;                                              // mm_interconnect_0:timer_2_s1_write -> timer_2:write_n
	wire  [15:0] mm_interconnect_0_timer_2_s1_writedata;                                          // mm_interconnect_0:timer_2_s1_writedata -> timer_2:writedata
	wire         mm_interconnect_0_esp32_spi_spi_control_port_chipselect;                         // mm_interconnect_0:esp32_spi_spi_control_port_chipselect -> esp32_spi:spi_select
	wire  [31:0] mm_interconnect_0_esp32_spi_spi_control_port_readdata;                           // esp32_spi:data_to_cpu -> mm_interconnect_0:esp32_spi_spi_control_port_readdata
	wire   [2:0] mm_interconnect_0_esp32_spi_spi_control_port_address;                            // mm_interconnect_0:esp32_spi_spi_control_port_address -> esp32_spi:mem_addr
	wire         mm_interconnect_0_esp32_spi_spi_control_port_read;                               // mm_interconnect_0:esp32_spi_spi_control_port_read -> esp32_spi:read_n
	wire         mm_interconnect_0_esp32_spi_spi_control_port_write;                              // mm_interconnect_0:esp32_spi_spi_control_port_write -> esp32_spi:write_n
	wire  [31:0] mm_interconnect_0_esp32_spi_spi_control_port_writedata;                          // mm_interconnect_0:esp32_spi_spi_control_port_writedata -> esp32_spi:data_from_cpu
	wire         irq_mapper_receiver0_irq;                                                        // accelerometer:irq -> irq_mapper:receiver0_irq
	wire         irq_mapper_receiver1_irq;                                                        // jtag:av_irq -> irq_mapper:receiver1_irq
	wire         irq_mapper_receiver2_irq;                                                        // esp32_spi:irq -> irq_mapper:receiver2_irq
	wire         irq_mapper_receiver3_irq;                                                        // sys_clk:irq -> irq_mapper:receiver3_irq
	wire         irq_mapper_receiver4_irq;                                                        // timer_1:irq -> irq_mapper:receiver4_irq
	wire         irq_mapper_receiver5_irq;                                                        // timer_2:irq -> irq_mapper:receiver5_irq
	wire  [31:0] nios2_cpu_irq_irq;                                                               // irq_mapper:sender_irq -> nios2_cpu:irq
	wire         rst_controller_reset_out_reset;                                                  // rst_controller:reset_out -> [accelerometer:reset, dram_controller:reset_n, esp32_spi:reset_n, irq_mapper:reset, jtag:rst_n, mm_interconnect_0:nios2_cpu_reset_reset_bridge_in_reset_reset, nios2_cpu:reset_n, rst_translator:in_reset, sys_clk:reset_n, timer_1:reset_n, timer_2:reset_n]
	wire         rst_controller_reset_out_reset_req;                                              // rst_controller:reset_req -> [nios2_cpu:reset_req, rst_translator:reset_req_in]
	wire         dram_clks_pll_reset_source_reset;                                                // dram_clks_pll:reset_source_reset -> rst_controller:reset_in0
	wire         rst_controller_001_reset_out_reset;                                              // rst_controller_001:reset_out -> dram_clks_pll:ref_reset_reset

	esp32SPIHardware_accelerometer accelerometer (
		.clk           (dram_clks_pll_sys_clk_clk),                                                       //                                 clk.clk
		.reset         (rst_controller_reset_out_reset),                                                  //                               reset.reset
		.address       (mm_interconnect_0_accelerometer_avalon_accelerometer_spi_mode_slave_address),     // avalon_accelerometer_spi_mode_slave.address
		.byteenable    (mm_interconnect_0_accelerometer_avalon_accelerometer_spi_mode_slave_byteenable),  //                                    .byteenable
		.read          (mm_interconnect_0_accelerometer_avalon_accelerometer_spi_mode_slave_read),        //                                    .read
		.write         (mm_interconnect_0_accelerometer_avalon_accelerometer_spi_mode_slave_write),       //                                    .write
		.writedata     (mm_interconnect_0_accelerometer_avalon_accelerometer_spi_mode_slave_writedata),   //                                    .writedata
		.readdata      (mm_interconnect_0_accelerometer_avalon_accelerometer_spi_mode_slave_readdata),    //                                    .readdata
		.waitrequest   (mm_interconnect_0_accelerometer_avalon_accelerometer_spi_mode_slave_waitrequest), //                                    .waitrequest
		.irq           (irq_mapper_receiver0_irq),                                                        //                           interrupt.irq
		.I2C_SDAT      (accelerometer_spi_I2C_SDAT),                                                      //                  external_interface.export
		.I2C_SCLK      (accelerometer_spi_I2C_SCLK),                                                      //                                    .export
		.G_SENSOR_CS_N (accelerometer_spi_G_SENSOR_CS_N),                                                 //                                    .export
		.G_SENSOR_INT  (accelerometer_spi_G_SENSOR_INT)                                                   //                                    .export
	);

	esp32SPIHardware_dram_clks_pll dram_clks_pll (
		.ref_clk_clk        (clk_clk),                            //      ref_clk.clk
		.ref_reset_reset    (rst_controller_001_reset_out_reset), //    ref_reset.reset
		.sys_clk_clk        (dram_clks_pll_sys_clk_clk),          //      sys_clk.clk
		.sdram_clk_clk      (sdram_clk_clk),                      //    sdram_clk.clk
		.reset_source_reset (dram_clks_pll_reset_source_reset)    // reset_source.reset
	);

	esp32SPIHardware_dram_controller dram_controller (
		.clk            (dram_clks_pll_sys_clk_clk),                          //   clk.clk
		.reset_n        (~rst_controller_reset_out_reset),                    // reset.reset_n
		.az_addr        (mm_interconnect_0_dram_controller_s1_address),       //    s1.address
		.az_be_n        (~mm_interconnect_0_dram_controller_s1_byteenable),   //      .byteenable_n
		.az_cs          (mm_interconnect_0_dram_controller_s1_chipselect),    //      .chipselect
		.az_data        (mm_interconnect_0_dram_controller_s1_writedata),     //      .writedata
		.az_rd_n        (~mm_interconnect_0_dram_controller_s1_read),         //      .read_n
		.az_wr_n        (~mm_interconnect_0_dram_controller_s1_write),        //      .write_n
		.za_data        (mm_interconnect_0_dram_controller_s1_readdata),      //      .readdata
		.za_valid       (mm_interconnect_0_dram_controller_s1_readdatavalid), //      .readdatavalid
		.za_waitrequest (mm_interconnect_0_dram_controller_s1_waitrequest),   //      .waitrequest
		.zs_addr        (dram_addr),                                          //  wire.export
		.zs_ba          (dram_ba),                                            //      .export
		.zs_cas_n       (dram_cas_n),                                         //      .export
		.zs_cke         (dram_cke),                                           //      .export
		.zs_cs_n        (dram_cs_n),                                          //      .export
		.zs_dq          (dram_dq),                                            //      .export
		.zs_dqm         (dram_dqm),                                           //      .export
		.zs_ras_n       (dram_ras_n),                                         //      .export
		.zs_we_n        (dram_we_n)                                           //      .export
	);

	esp32SPIHardware_esp32_spi esp32_spi (
		.clk           (dram_clks_pll_sys_clk_clk),                               //              clk.clk
		.reset_n       (~rst_controller_reset_out_reset),                         //            reset.reset_n
		.data_from_cpu (mm_interconnect_0_esp32_spi_spi_control_port_writedata),  // spi_control_port.writedata
		.data_to_cpu   (mm_interconnect_0_esp32_spi_spi_control_port_readdata),   //                 .readdata
		.mem_addr      (mm_interconnect_0_esp32_spi_spi_control_port_address),    //                 .address
		.read_n        (~mm_interconnect_0_esp32_spi_spi_control_port_read),      //                 .read_n
		.spi_select    (mm_interconnect_0_esp32_spi_spi_control_port_chipselect), //                 .chipselect
		.write_n       (~mm_interconnect_0_esp32_spi_spi_control_port_write),     //                 .write_n
		.irq           (irq_mapper_receiver2_irq),                                //              irq.irq
		.MISO          (esp32_spi_MISO),                                          //         external.export
		.MOSI          (esp32_spi_MOSI),                                          //                 .export
		.SCLK          (esp32_spi_SCLK),                                          //                 .export
		.SS_n          (esp32_spi_SS_n)                                           //                 .export
	);

	esp32SPIHardware_fph2 #(
		.arithmetic_present (1),
		.root_present       (0),
		.conversion_present (1),
		.comparison_present (1)
	) fph2 (
		.s1_dataa     (nios2_cpu_custom_instruction_master_comb_slave_translator0_ci_master_dataa),      // s1.dataa
		.s1_datab     (nios2_cpu_custom_instruction_master_comb_slave_translator0_ci_master_datab),      //   .datab
		.s1_n         (nios2_cpu_custom_instruction_master_comb_slave_translator0_ci_master_n),          //   .n
		.s1_result    (nios2_cpu_custom_instruction_master_comb_slave_translator0_ci_master_result),     //   .result
		.s2_clk       (nios2_cpu_custom_instruction_master_multi_slave_translator0_ci_master_clk),       // s2.clk
		.s2_clk_en    (nios2_cpu_custom_instruction_master_multi_slave_translator0_ci_master_clk_en),    //   .clk_en
		.s2_dataa     (nios2_cpu_custom_instruction_master_multi_slave_translator0_ci_master_dataa),     //   .dataa
		.s2_datab     (nios2_cpu_custom_instruction_master_multi_slave_translator0_ci_master_datab),     //   .datab
		.s2_n         (nios2_cpu_custom_instruction_master_multi_slave_translator0_ci_master_n),         //   .n
		.s2_reset     (nios2_cpu_custom_instruction_master_multi_slave_translator0_ci_master_reset),     //   .reset
		.s2_reset_req (nios2_cpu_custom_instruction_master_multi_slave_translator0_ci_master_reset_req), //   .reset_req
		.s2_start     (nios2_cpu_custom_instruction_master_multi_slave_translator0_ci_master_start),     //   .start
		.s2_done      (nios2_cpu_custom_instruction_master_multi_slave_translator0_ci_master_done),      //   .done
		.s2_result    (nios2_cpu_custom_instruction_master_multi_slave_translator0_ci_master_result)     //   .result
	);

	esp32SPIHardware_jtag jtag (
		.clk            (dram_clks_pll_sys_clk_clk),                            //               clk.clk
		.rst_n          (~rst_controller_reset_out_reset),                      //             reset.reset_n
		.av_chipselect  (mm_interconnect_0_jtag_avalon_jtag_slave_chipselect),  // avalon_jtag_slave.chipselect
		.av_address     (mm_interconnect_0_jtag_avalon_jtag_slave_address),     //                  .address
		.av_read_n      (~mm_interconnect_0_jtag_avalon_jtag_slave_read),       //                  .read_n
		.av_readdata    (mm_interconnect_0_jtag_avalon_jtag_slave_readdata),    //                  .readdata
		.av_write_n     (~mm_interconnect_0_jtag_avalon_jtag_slave_write),      //                  .write_n
		.av_writedata   (mm_interconnect_0_jtag_avalon_jtag_slave_writedata),   //                  .writedata
		.av_waitrequest (mm_interconnect_0_jtag_avalon_jtag_slave_waitrequest), //                  .waitrequest
		.av_irq         (irq_mapper_receiver1_irq)                              //               irq.irq
	);

	esp32SPIHardware_nios2_cpu nios2_cpu (
		.clk                                 (dram_clks_pll_sys_clk_clk),                               //                       clk.clk
		.reset_n                             (~rst_controller_reset_out_reset),                         //                     reset.reset_n
		.reset_req                           (rst_controller_reset_out_reset_req),                      //                          .reset_req
		.d_address                           (nios2_cpu_data_master_address),                           //               data_master.address
		.d_byteenable                        (nios2_cpu_data_master_byteenable),                        //                          .byteenable
		.d_read                              (nios2_cpu_data_master_read),                              //                          .read
		.d_readdata                          (nios2_cpu_data_master_readdata),                          //                          .readdata
		.d_waitrequest                       (nios2_cpu_data_master_waitrequest),                       //                          .waitrequest
		.d_write                             (nios2_cpu_data_master_write),                             //                          .write
		.d_writedata                         (nios2_cpu_data_master_writedata),                         //                          .writedata
		.d_readdatavalid                     (nios2_cpu_data_master_readdatavalid),                     //                          .readdatavalid
		.debug_mem_slave_debugaccess_to_roms (nios2_cpu_data_master_debugaccess),                       //                          .debugaccess
		.i_address                           (nios2_cpu_instruction_master_address),                    //        instruction_master.address
		.i_read                              (nios2_cpu_instruction_master_read),                       //                          .read
		.i_readdata                          (nios2_cpu_instruction_master_readdata),                   //                          .readdata
		.i_waitrequest                       (nios2_cpu_instruction_master_waitrequest),                //                          .waitrequest
		.i_readdatavalid                     (nios2_cpu_instruction_master_readdatavalid),              //                          .readdatavalid
		.irq                                 (nios2_cpu_irq_irq),                                       //                       irq.irq
		.debug_reset_request                 (),                                                        //       debug_reset_request.reset
		.debug_mem_slave_address             (mm_interconnect_0_nios2_cpu_debug_mem_slave_address),     //           debug_mem_slave.address
		.debug_mem_slave_byteenable          (mm_interconnect_0_nios2_cpu_debug_mem_slave_byteenable),  //                          .byteenable
		.debug_mem_slave_debugaccess         (mm_interconnect_0_nios2_cpu_debug_mem_slave_debugaccess), //                          .debugaccess
		.debug_mem_slave_read                (mm_interconnect_0_nios2_cpu_debug_mem_slave_read),        //                          .read
		.debug_mem_slave_readdata            (mm_interconnect_0_nios2_cpu_debug_mem_slave_readdata),    //                          .readdata
		.debug_mem_slave_waitrequest         (mm_interconnect_0_nios2_cpu_debug_mem_slave_waitrequest), //                          .waitrequest
		.debug_mem_slave_write               (mm_interconnect_0_nios2_cpu_debug_mem_slave_write),       //                          .write
		.debug_mem_slave_writedata           (mm_interconnect_0_nios2_cpu_debug_mem_slave_writedata),   //                          .writedata
		.A_ci_multi_done                     (nios2_cpu_custom_instruction_master_done),                // custom_instruction_master.done
		.A_ci_multi_result                   (nios2_cpu_custom_instruction_master_multi_result),        //                          .multi_result
		.A_ci_multi_a                        (nios2_cpu_custom_instruction_master_multi_a),             //                          .multi_a
		.A_ci_multi_b                        (nios2_cpu_custom_instruction_master_multi_b),             //                          .multi_b
		.A_ci_multi_c                        (nios2_cpu_custom_instruction_master_multi_c),             //                          .multi_c
		.A_ci_multi_clk_en                   (nios2_cpu_custom_instruction_master_clk_en),              //                          .clk_en
		.A_ci_multi_clock                    (nios2_cpu_custom_instruction_master_clk),                 //                          .clk
		.A_ci_multi_reset                    (nios2_cpu_custom_instruction_master_reset),               //                          .reset
		.A_ci_multi_reset_req                (nios2_cpu_custom_instruction_master_reset_req),           //                          .reset_req
		.A_ci_multi_dataa                    (nios2_cpu_custom_instruction_master_multi_dataa),         //                          .multi_dataa
		.A_ci_multi_datab                    (nios2_cpu_custom_instruction_master_multi_datab),         //                          .multi_datab
		.A_ci_multi_n                        (nios2_cpu_custom_instruction_master_multi_n),             //                          .multi_n
		.A_ci_multi_readra                   (nios2_cpu_custom_instruction_master_multi_readra),        //                          .multi_readra
		.A_ci_multi_readrb                   (nios2_cpu_custom_instruction_master_multi_readrb),        //                          .multi_readrb
		.A_ci_multi_start                    (nios2_cpu_custom_instruction_master_start),               //                          .start
		.A_ci_multi_writerc                  (nios2_cpu_custom_instruction_master_multi_writerc),       //                          .multi_writerc
		.E_ci_combo_result                   (nios2_cpu_custom_instruction_master_result),              //                          .result
		.E_ci_combo_a                        (nios2_cpu_custom_instruction_master_a),                   //                          .a
		.E_ci_combo_b                        (nios2_cpu_custom_instruction_master_b),                   //                          .b
		.E_ci_combo_c                        (nios2_cpu_custom_instruction_master_c),                   //                          .c
		.E_ci_combo_dataa                    (nios2_cpu_custom_instruction_master_dataa),               //                          .dataa
		.E_ci_combo_datab                    (nios2_cpu_custom_instruction_master_datab),               //                          .datab
		.E_ci_combo_estatus                  (nios2_cpu_custom_instruction_master_estatus),             //                          .estatus
		.E_ci_combo_ipending                 (nios2_cpu_custom_instruction_master_ipending),            //                          .ipending
		.E_ci_combo_n                        (nios2_cpu_custom_instruction_master_n),                   //                          .n
		.E_ci_combo_readra                   (nios2_cpu_custom_instruction_master_readra),              //                          .readra
		.E_ci_combo_readrb                   (nios2_cpu_custom_instruction_master_readrb),              //                          .readrb
		.E_ci_combo_writerc                  (nios2_cpu_custom_instruction_master_writerc)              //                          .writerc
	);

	esp32SPIHardware_sys_clk sys_clk (
		.clk        (dram_clks_pll_sys_clk_clk),               //   clk.clk
		.reset_n    (~rst_controller_reset_out_reset),         // reset.reset_n
		.address    (mm_interconnect_0_sys_clk_s1_address),    //    s1.address
		.writedata  (mm_interconnect_0_sys_clk_s1_writedata),  //      .writedata
		.readdata   (mm_interconnect_0_sys_clk_s1_readdata),   //      .readdata
		.chipselect (mm_interconnect_0_sys_clk_s1_chipselect), //      .chipselect
		.write_n    (~mm_interconnect_0_sys_clk_s1_write),     //      .write_n
		.irq        (irq_mapper_receiver3_irq)                 //   irq.irq
	);

	esp32SPIHardware_sys_clk timer_1 (
		.clk        (dram_clks_pll_sys_clk_clk),               //   clk.clk
		.reset_n    (~rst_controller_reset_out_reset),         // reset.reset_n
		.address    (mm_interconnect_0_timer_1_s1_address),    //    s1.address
		.writedata  (mm_interconnect_0_timer_1_s1_writedata),  //      .writedata
		.readdata   (mm_interconnect_0_timer_1_s1_readdata),   //      .readdata
		.chipselect (mm_interconnect_0_timer_1_s1_chipselect), //      .chipselect
		.write_n    (~mm_interconnect_0_timer_1_s1_write),     //      .write_n
		.irq        (irq_mapper_receiver4_irq)                 //   irq.irq
	);

	esp32SPIHardware_sys_clk timer_2 (
		.clk        (dram_clks_pll_sys_clk_clk),               //   clk.clk
		.reset_n    (~rst_controller_reset_out_reset),         // reset.reset_n
		.address    (mm_interconnect_0_timer_2_s1_address),    //    s1.address
		.writedata  (mm_interconnect_0_timer_2_s1_writedata),  //      .writedata
		.readdata   (mm_interconnect_0_timer_2_s1_readdata),   //      .readdata
		.chipselect (mm_interconnect_0_timer_2_s1_chipselect), //      .chipselect
		.write_n    (~mm_interconnect_0_timer_2_s1_write),     //      .write_n
		.irq        (irq_mapper_receiver5_irq)                 //   irq.irq
	);

	altera_customins_master_translator #(
		.SHARED_COMB_AND_MULTI (0)
	) nios2_cpu_custom_instruction_master_translator (
		.ci_slave_dataa            (nios2_cpu_custom_instruction_master_dataa),                                //        ci_slave.dataa
		.ci_slave_datab            (nios2_cpu_custom_instruction_master_datab),                                //                .datab
		.ci_slave_result           (nios2_cpu_custom_instruction_master_result),                               //                .result
		.ci_slave_n                (nios2_cpu_custom_instruction_master_n),                                    //                .n
		.ci_slave_readra           (nios2_cpu_custom_instruction_master_readra),                               //                .readra
		.ci_slave_readrb           (nios2_cpu_custom_instruction_master_readrb),                               //                .readrb
		.ci_slave_writerc          (nios2_cpu_custom_instruction_master_writerc),                              //                .writerc
		.ci_slave_a                (nios2_cpu_custom_instruction_master_a),                                    //                .a
		.ci_slave_b                (nios2_cpu_custom_instruction_master_b),                                    //                .b
		.ci_slave_c                (nios2_cpu_custom_instruction_master_c),                                    //                .c
		.ci_slave_ipending         (nios2_cpu_custom_instruction_master_ipending),                             //                .ipending
		.ci_slave_estatus          (nios2_cpu_custom_instruction_master_estatus),                              //                .estatus
		.ci_slave_multi_clk        (nios2_cpu_custom_instruction_master_clk),                                  //                .clk
		.ci_slave_multi_reset      (nios2_cpu_custom_instruction_master_reset),                                //                .reset
		.ci_slave_multi_clken      (nios2_cpu_custom_instruction_master_clk_en),                               //                .clk_en
		.ci_slave_multi_reset_req  (nios2_cpu_custom_instruction_master_reset_req),                            //                .reset_req
		.ci_slave_multi_start      (nios2_cpu_custom_instruction_master_start),                                //                .start
		.ci_slave_multi_done       (nios2_cpu_custom_instruction_master_done),                                 //                .done
		.ci_slave_multi_dataa      (nios2_cpu_custom_instruction_master_multi_dataa),                          //                .multi_dataa
		.ci_slave_multi_datab      (nios2_cpu_custom_instruction_master_multi_datab),                          //                .multi_datab
		.ci_slave_multi_result     (nios2_cpu_custom_instruction_master_multi_result),                         //                .multi_result
		.ci_slave_multi_n          (nios2_cpu_custom_instruction_master_multi_n),                              //                .multi_n
		.ci_slave_multi_readra     (nios2_cpu_custom_instruction_master_multi_readra),                         //                .multi_readra
		.ci_slave_multi_readrb     (nios2_cpu_custom_instruction_master_multi_readrb),                         //                .multi_readrb
		.ci_slave_multi_writerc    (nios2_cpu_custom_instruction_master_multi_writerc),                        //                .multi_writerc
		.ci_slave_multi_a          (nios2_cpu_custom_instruction_master_multi_a),                              //                .multi_a
		.ci_slave_multi_b          (nios2_cpu_custom_instruction_master_multi_b),                              //                .multi_b
		.ci_slave_multi_c          (nios2_cpu_custom_instruction_master_multi_c),                              //                .multi_c
		.comb_ci_master_dataa      (nios2_cpu_custom_instruction_master_translator_comb_ci_master_dataa),      //  comb_ci_master.dataa
		.comb_ci_master_datab      (nios2_cpu_custom_instruction_master_translator_comb_ci_master_datab),      //                .datab
		.comb_ci_master_result     (nios2_cpu_custom_instruction_master_translator_comb_ci_master_result),     //                .result
		.comb_ci_master_n          (nios2_cpu_custom_instruction_master_translator_comb_ci_master_n),          //                .n
		.comb_ci_master_readra     (nios2_cpu_custom_instruction_master_translator_comb_ci_master_readra),     //                .readra
		.comb_ci_master_readrb     (nios2_cpu_custom_instruction_master_translator_comb_ci_master_readrb),     //                .readrb
		.comb_ci_master_writerc    (nios2_cpu_custom_instruction_master_translator_comb_ci_master_writerc),    //                .writerc
		.comb_ci_master_a          (nios2_cpu_custom_instruction_master_translator_comb_ci_master_a),          //                .a
		.comb_ci_master_b          (nios2_cpu_custom_instruction_master_translator_comb_ci_master_b),          //                .b
		.comb_ci_master_c          (nios2_cpu_custom_instruction_master_translator_comb_ci_master_c),          //                .c
		.comb_ci_master_ipending   (nios2_cpu_custom_instruction_master_translator_comb_ci_master_ipending),   //                .ipending
		.comb_ci_master_estatus    (nios2_cpu_custom_instruction_master_translator_comb_ci_master_estatus),    //                .estatus
		.multi_ci_master_clk       (nios2_cpu_custom_instruction_master_translator_multi_ci_master_clk),       // multi_ci_master.clk
		.multi_ci_master_reset     (nios2_cpu_custom_instruction_master_translator_multi_ci_master_reset),     //                .reset
		.multi_ci_master_clken     (nios2_cpu_custom_instruction_master_translator_multi_ci_master_clk_en),    //                .clk_en
		.multi_ci_master_reset_req (nios2_cpu_custom_instruction_master_translator_multi_ci_master_reset_req), //                .reset_req
		.multi_ci_master_start     (nios2_cpu_custom_instruction_master_translator_multi_ci_master_start),     //                .start
		.multi_ci_master_done      (nios2_cpu_custom_instruction_master_translator_multi_ci_master_done),      //                .done
		.multi_ci_master_dataa     (nios2_cpu_custom_instruction_master_translator_multi_ci_master_dataa),     //                .dataa
		.multi_ci_master_datab     (nios2_cpu_custom_instruction_master_translator_multi_ci_master_datab),     //                .datab
		.multi_ci_master_result    (nios2_cpu_custom_instruction_master_translator_multi_ci_master_result),    //                .result
		.multi_ci_master_n         (nios2_cpu_custom_instruction_master_translator_multi_ci_master_n),         //                .n
		.multi_ci_master_readra    (nios2_cpu_custom_instruction_master_translator_multi_ci_master_readra),    //                .readra
		.multi_ci_master_readrb    (nios2_cpu_custom_instruction_master_translator_multi_ci_master_readrb),    //                .readrb
		.multi_ci_master_writerc   (nios2_cpu_custom_instruction_master_translator_multi_ci_master_writerc),   //                .writerc
		.multi_ci_master_a         (nios2_cpu_custom_instruction_master_translator_multi_ci_master_a),         //                .a
		.multi_ci_master_b         (nios2_cpu_custom_instruction_master_translator_multi_ci_master_b),         //                .b
		.multi_ci_master_c         (nios2_cpu_custom_instruction_master_translator_multi_ci_master_c)          //                .c
	);

	esp32SPIHardware_nios2_cpu_custom_instruction_master_comb_xconnect nios2_cpu_custom_instruction_master_comb_xconnect (
		.ci_slave_dataa      (nios2_cpu_custom_instruction_master_translator_comb_ci_master_dataa),    //   ci_slave.dataa
		.ci_slave_datab      (nios2_cpu_custom_instruction_master_translator_comb_ci_master_datab),    //           .datab
		.ci_slave_result     (nios2_cpu_custom_instruction_master_translator_comb_ci_master_result),   //           .result
		.ci_slave_n          (nios2_cpu_custom_instruction_master_translator_comb_ci_master_n),        //           .n
		.ci_slave_readra     (nios2_cpu_custom_instruction_master_translator_comb_ci_master_readra),   //           .readra
		.ci_slave_readrb     (nios2_cpu_custom_instruction_master_translator_comb_ci_master_readrb),   //           .readrb
		.ci_slave_writerc    (nios2_cpu_custom_instruction_master_translator_comb_ci_master_writerc),  //           .writerc
		.ci_slave_a          (nios2_cpu_custom_instruction_master_translator_comb_ci_master_a),        //           .a
		.ci_slave_b          (nios2_cpu_custom_instruction_master_translator_comb_ci_master_b),        //           .b
		.ci_slave_c          (nios2_cpu_custom_instruction_master_translator_comb_ci_master_c),        //           .c
		.ci_slave_ipending   (nios2_cpu_custom_instruction_master_translator_comb_ci_master_ipending), //           .ipending
		.ci_slave_estatus    (nios2_cpu_custom_instruction_master_translator_comb_ci_master_estatus),  //           .estatus
		.ci_master0_dataa    (nios2_cpu_custom_instruction_master_comb_xconnect_ci_master0_dataa),     // ci_master0.dataa
		.ci_master0_datab    (nios2_cpu_custom_instruction_master_comb_xconnect_ci_master0_datab),     //           .datab
		.ci_master0_result   (nios2_cpu_custom_instruction_master_comb_xconnect_ci_master0_result),    //           .result
		.ci_master0_n        (nios2_cpu_custom_instruction_master_comb_xconnect_ci_master0_n),         //           .n
		.ci_master0_readra   (nios2_cpu_custom_instruction_master_comb_xconnect_ci_master0_readra),    //           .readra
		.ci_master0_readrb   (nios2_cpu_custom_instruction_master_comb_xconnect_ci_master0_readrb),    //           .readrb
		.ci_master0_writerc  (nios2_cpu_custom_instruction_master_comb_xconnect_ci_master0_writerc),   //           .writerc
		.ci_master0_a        (nios2_cpu_custom_instruction_master_comb_xconnect_ci_master0_a),         //           .a
		.ci_master0_b        (nios2_cpu_custom_instruction_master_comb_xconnect_ci_master0_b),         //           .b
		.ci_master0_c        (nios2_cpu_custom_instruction_master_comb_xconnect_ci_master0_c),         //           .c
		.ci_master0_ipending (nios2_cpu_custom_instruction_master_comb_xconnect_ci_master0_ipending),  //           .ipending
		.ci_master0_estatus  (nios2_cpu_custom_instruction_master_comb_xconnect_ci_master0_estatus)    //           .estatus
	);

	altera_customins_slave_translator #(
		.N_WIDTH          (4),
		.USE_DONE         (0),
		.NUM_FIXED_CYCLES (0)
	) nios2_cpu_custom_instruction_master_comb_slave_translator0 (
		.ci_slave_dataa      (nios2_cpu_custom_instruction_master_comb_xconnect_ci_master0_dataa),          //  ci_slave.dataa
		.ci_slave_datab      (nios2_cpu_custom_instruction_master_comb_xconnect_ci_master0_datab),          //          .datab
		.ci_slave_result     (nios2_cpu_custom_instruction_master_comb_xconnect_ci_master0_result),         //          .result
		.ci_slave_n          (nios2_cpu_custom_instruction_master_comb_xconnect_ci_master0_n),              //          .n
		.ci_slave_readra     (nios2_cpu_custom_instruction_master_comb_xconnect_ci_master0_readra),         //          .readra
		.ci_slave_readrb     (nios2_cpu_custom_instruction_master_comb_xconnect_ci_master0_readrb),         //          .readrb
		.ci_slave_writerc    (nios2_cpu_custom_instruction_master_comb_xconnect_ci_master0_writerc),        //          .writerc
		.ci_slave_a          (nios2_cpu_custom_instruction_master_comb_xconnect_ci_master0_a),              //          .a
		.ci_slave_b          (nios2_cpu_custom_instruction_master_comb_xconnect_ci_master0_b),              //          .b
		.ci_slave_c          (nios2_cpu_custom_instruction_master_comb_xconnect_ci_master0_c),              //          .c
		.ci_slave_ipending   (nios2_cpu_custom_instruction_master_comb_xconnect_ci_master0_ipending),       //          .ipending
		.ci_slave_estatus    (nios2_cpu_custom_instruction_master_comb_xconnect_ci_master0_estatus),        //          .estatus
		.ci_master_dataa     (nios2_cpu_custom_instruction_master_comb_slave_translator0_ci_master_dataa),  // ci_master.dataa
		.ci_master_datab     (nios2_cpu_custom_instruction_master_comb_slave_translator0_ci_master_datab),  //          .datab
		.ci_master_result    (nios2_cpu_custom_instruction_master_comb_slave_translator0_ci_master_result), //          .result
		.ci_master_n         (nios2_cpu_custom_instruction_master_comb_slave_translator0_ci_master_n),      //          .n
		.ci_master_readra    (),                                                                            // (terminated)
		.ci_master_readrb    (),                                                                            // (terminated)
		.ci_master_writerc   (),                                                                            // (terminated)
		.ci_master_a         (),                                                                            // (terminated)
		.ci_master_b         (),                                                                            // (terminated)
		.ci_master_c         (),                                                                            // (terminated)
		.ci_master_ipending  (),                                                                            // (terminated)
		.ci_master_estatus   (),                                                                            // (terminated)
		.ci_master_clk       (),                                                                            // (terminated)
		.ci_master_clken     (),                                                                            // (terminated)
		.ci_master_reset_req (),                                                                            // (terminated)
		.ci_master_reset     (),                                                                            // (terminated)
		.ci_master_start     (),                                                                            // (terminated)
		.ci_master_done      (1'b0),                                                                        // (terminated)
		.ci_slave_clk        (1'b0),                                                                        // (terminated)
		.ci_slave_clken      (1'b0),                                                                        // (terminated)
		.ci_slave_reset_req  (1'b0),                                                                        // (terminated)
		.ci_slave_reset      (1'b0),                                                                        // (terminated)
		.ci_slave_start      (1'b0),                                                                        // (terminated)
		.ci_slave_done       ()                                                                             // (terminated)
	);

	esp32SPIHardware_nios2_cpu_custom_instruction_master_multi_xconnect nios2_cpu_custom_instruction_master_multi_xconnect (
		.ci_slave_dataa       (nios2_cpu_custom_instruction_master_translator_multi_ci_master_dataa),     //   ci_slave.dataa
		.ci_slave_datab       (nios2_cpu_custom_instruction_master_translator_multi_ci_master_datab),     //           .datab
		.ci_slave_result      (nios2_cpu_custom_instruction_master_translator_multi_ci_master_result),    //           .result
		.ci_slave_n           (nios2_cpu_custom_instruction_master_translator_multi_ci_master_n),         //           .n
		.ci_slave_readra      (nios2_cpu_custom_instruction_master_translator_multi_ci_master_readra),    //           .readra
		.ci_slave_readrb      (nios2_cpu_custom_instruction_master_translator_multi_ci_master_readrb),    //           .readrb
		.ci_slave_writerc     (nios2_cpu_custom_instruction_master_translator_multi_ci_master_writerc),   //           .writerc
		.ci_slave_a           (nios2_cpu_custom_instruction_master_translator_multi_ci_master_a),         //           .a
		.ci_slave_b           (nios2_cpu_custom_instruction_master_translator_multi_ci_master_b),         //           .b
		.ci_slave_c           (nios2_cpu_custom_instruction_master_translator_multi_ci_master_c),         //           .c
		.ci_slave_ipending    (),                                                                         //           .ipending
		.ci_slave_estatus     (),                                                                         //           .estatus
		.ci_slave_clk         (nios2_cpu_custom_instruction_master_translator_multi_ci_master_clk),       //           .clk
		.ci_slave_reset       (nios2_cpu_custom_instruction_master_translator_multi_ci_master_reset),     //           .reset
		.ci_slave_clken       (nios2_cpu_custom_instruction_master_translator_multi_ci_master_clk_en),    //           .clk_en
		.ci_slave_reset_req   (nios2_cpu_custom_instruction_master_translator_multi_ci_master_reset_req), //           .reset_req
		.ci_slave_start       (nios2_cpu_custom_instruction_master_translator_multi_ci_master_start),     //           .start
		.ci_slave_done        (nios2_cpu_custom_instruction_master_translator_multi_ci_master_done),      //           .done
		.ci_master0_dataa     (nios2_cpu_custom_instruction_master_multi_xconnect_ci_master0_dataa),      // ci_master0.dataa
		.ci_master0_datab     (nios2_cpu_custom_instruction_master_multi_xconnect_ci_master0_datab),      //           .datab
		.ci_master0_result    (nios2_cpu_custom_instruction_master_multi_xconnect_ci_master0_result),     //           .result
		.ci_master0_n         (nios2_cpu_custom_instruction_master_multi_xconnect_ci_master0_n),          //           .n
		.ci_master0_readra    (nios2_cpu_custom_instruction_master_multi_xconnect_ci_master0_readra),     //           .readra
		.ci_master0_readrb    (nios2_cpu_custom_instruction_master_multi_xconnect_ci_master0_readrb),     //           .readrb
		.ci_master0_writerc   (nios2_cpu_custom_instruction_master_multi_xconnect_ci_master0_writerc),    //           .writerc
		.ci_master0_a         (nios2_cpu_custom_instruction_master_multi_xconnect_ci_master0_a),          //           .a
		.ci_master0_b         (nios2_cpu_custom_instruction_master_multi_xconnect_ci_master0_b),          //           .b
		.ci_master0_c         (nios2_cpu_custom_instruction_master_multi_xconnect_ci_master0_c),          //           .c
		.ci_master0_ipending  (nios2_cpu_custom_instruction_master_multi_xconnect_ci_master0_ipending),   //           .ipending
		.ci_master0_estatus   (nios2_cpu_custom_instruction_master_multi_xconnect_ci_master0_estatus),    //           .estatus
		.ci_master0_clk       (nios2_cpu_custom_instruction_master_multi_xconnect_ci_master0_clk),        //           .clk
		.ci_master0_reset     (nios2_cpu_custom_instruction_master_multi_xconnect_ci_master0_reset),      //           .reset
		.ci_master0_clken     (nios2_cpu_custom_instruction_master_multi_xconnect_ci_master0_clk_en),     //           .clk_en
		.ci_master0_reset_req (nios2_cpu_custom_instruction_master_multi_xconnect_ci_master0_reset_req),  //           .reset_req
		.ci_master0_start     (nios2_cpu_custom_instruction_master_multi_xconnect_ci_master0_start),      //           .start
		.ci_master0_done      (nios2_cpu_custom_instruction_master_multi_xconnect_ci_master0_done)        //           .done
	);

	altera_customins_slave_translator #(
		.N_WIDTH          (3),
		.USE_DONE         (1),
		.NUM_FIXED_CYCLES (1)
	) nios2_cpu_custom_instruction_master_multi_slave_translator0 (
		.ci_slave_dataa      (nios2_cpu_custom_instruction_master_multi_xconnect_ci_master0_dataa),             //  ci_slave.dataa
		.ci_slave_datab      (nios2_cpu_custom_instruction_master_multi_xconnect_ci_master0_datab),             //          .datab
		.ci_slave_result     (nios2_cpu_custom_instruction_master_multi_xconnect_ci_master0_result),            //          .result
		.ci_slave_n          (nios2_cpu_custom_instruction_master_multi_xconnect_ci_master0_n),                 //          .n
		.ci_slave_readra     (nios2_cpu_custom_instruction_master_multi_xconnect_ci_master0_readra),            //          .readra
		.ci_slave_readrb     (nios2_cpu_custom_instruction_master_multi_xconnect_ci_master0_readrb),            //          .readrb
		.ci_slave_writerc    (nios2_cpu_custom_instruction_master_multi_xconnect_ci_master0_writerc),           //          .writerc
		.ci_slave_a          (nios2_cpu_custom_instruction_master_multi_xconnect_ci_master0_a),                 //          .a
		.ci_slave_b          (nios2_cpu_custom_instruction_master_multi_xconnect_ci_master0_b),                 //          .b
		.ci_slave_c          (nios2_cpu_custom_instruction_master_multi_xconnect_ci_master0_c),                 //          .c
		.ci_slave_ipending   (nios2_cpu_custom_instruction_master_multi_xconnect_ci_master0_ipending),          //          .ipending
		.ci_slave_estatus    (nios2_cpu_custom_instruction_master_multi_xconnect_ci_master0_estatus),           //          .estatus
		.ci_slave_clk        (nios2_cpu_custom_instruction_master_multi_xconnect_ci_master0_clk),               //          .clk
		.ci_slave_clken      (nios2_cpu_custom_instruction_master_multi_xconnect_ci_master0_clk_en),            //          .clk_en
		.ci_slave_reset_req  (nios2_cpu_custom_instruction_master_multi_xconnect_ci_master0_reset_req),         //          .reset_req
		.ci_slave_reset      (nios2_cpu_custom_instruction_master_multi_xconnect_ci_master0_reset),             //          .reset
		.ci_slave_start      (nios2_cpu_custom_instruction_master_multi_xconnect_ci_master0_start),             //          .start
		.ci_slave_done       (nios2_cpu_custom_instruction_master_multi_xconnect_ci_master0_done),              //          .done
		.ci_master_dataa     (nios2_cpu_custom_instruction_master_multi_slave_translator0_ci_master_dataa),     // ci_master.dataa
		.ci_master_datab     (nios2_cpu_custom_instruction_master_multi_slave_translator0_ci_master_datab),     //          .datab
		.ci_master_result    (nios2_cpu_custom_instruction_master_multi_slave_translator0_ci_master_result),    //          .result
		.ci_master_n         (nios2_cpu_custom_instruction_master_multi_slave_translator0_ci_master_n),         //          .n
		.ci_master_clk       (nios2_cpu_custom_instruction_master_multi_slave_translator0_ci_master_clk),       //          .clk
		.ci_master_clken     (nios2_cpu_custom_instruction_master_multi_slave_translator0_ci_master_clk_en),    //          .clk_en
		.ci_master_reset_req (nios2_cpu_custom_instruction_master_multi_slave_translator0_ci_master_reset_req), //          .reset_req
		.ci_master_reset     (nios2_cpu_custom_instruction_master_multi_slave_translator0_ci_master_reset),     //          .reset
		.ci_master_start     (nios2_cpu_custom_instruction_master_multi_slave_translator0_ci_master_start),     //          .start
		.ci_master_done      (nios2_cpu_custom_instruction_master_multi_slave_translator0_ci_master_done),      //          .done
		.ci_master_readra    (),                                                                                // (terminated)
		.ci_master_readrb    (),                                                                                // (terminated)
		.ci_master_writerc   (),                                                                                // (terminated)
		.ci_master_a         (),                                                                                // (terminated)
		.ci_master_b         (),                                                                                // (terminated)
		.ci_master_c         (),                                                                                // (terminated)
		.ci_master_ipending  (),                                                                                // (terminated)
		.ci_master_estatus   ()                                                                                 // (terminated)
	);

	esp32SPIHardware_mm_interconnect_0 mm_interconnect_0 (
		.dram_clks_pll_sys_clk_clk                                     (dram_clks_pll_sys_clk_clk),                                                       //                             dram_clks_pll_sys_clk.clk
		.nios2_cpu_reset_reset_bridge_in_reset_reset                   (rst_controller_reset_out_reset),                                                  //             nios2_cpu_reset_reset_bridge_in_reset.reset
		.nios2_cpu_data_master_address                                 (nios2_cpu_data_master_address),                                                   //                             nios2_cpu_data_master.address
		.nios2_cpu_data_master_waitrequest                             (nios2_cpu_data_master_waitrequest),                                               //                                                  .waitrequest
		.nios2_cpu_data_master_byteenable                              (nios2_cpu_data_master_byteenable),                                                //                                                  .byteenable
		.nios2_cpu_data_master_read                                    (nios2_cpu_data_master_read),                                                      //                                                  .read
		.nios2_cpu_data_master_readdata                                (nios2_cpu_data_master_readdata),                                                  //                                                  .readdata
		.nios2_cpu_data_master_readdatavalid                           (nios2_cpu_data_master_readdatavalid),                                             //                                                  .readdatavalid
		.nios2_cpu_data_master_write                                   (nios2_cpu_data_master_write),                                                     //                                                  .write
		.nios2_cpu_data_master_writedata                               (nios2_cpu_data_master_writedata),                                                 //                                                  .writedata
		.nios2_cpu_data_master_debugaccess                             (nios2_cpu_data_master_debugaccess),                                               //                                                  .debugaccess
		.nios2_cpu_instruction_master_address                          (nios2_cpu_instruction_master_address),                                            //                      nios2_cpu_instruction_master.address
		.nios2_cpu_instruction_master_waitrequest                      (nios2_cpu_instruction_master_waitrequest),                                        //                                                  .waitrequest
		.nios2_cpu_instruction_master_read                             (nios2_cpu_instruction_master_read),                                               //                                                  .read
		.nios2_cpu_instruction_master_readdata                         (nios2_cpu_instruction_master_readdata),                                           //                                                  .readdata
		.nios2_cpu_instruction_master_readdatavalid                    (nios2_cpu_instruction_master_readdatavalid),                                      //                                                  .readdatavalid
		.accelerometer_avalon_accelerometer_spi_mode_slave_address     (mm_interconnect_0_accelerometer_avalon_accelerometer_spi_mode_slave_address),     // accelerometer_avalon_accelerometer_spi_mode_slave.address
		.accelerometer_avalon_accelerometer_spi_mode_slave_write       (mm_interconnect_0_accelerometer_avalon_accelerometer_spi_mode_slave_write),       //                                                  .write
		.accelerometer_avalon_accelerometer_spi_mode_slave_read        (mm_interconnect_0_accelerometer_avalon_accelerometer_spi_mode_slave_read),        //                                                  .read
		.accelerometer_avalon_accelerometer_spi_mode_slave_readdata    (mm_interconnect_0_accelerometer_avalon_accelerometer_spi_mode_slave_readdata),    //                                                  .readdata
		.accelerometer_avalon_accelerometer_spi_mode_slave_writedata   (mm_interconnect_0_accelerometer_avalon_accelerometer_spi_mode_slave_writedata),   //                                                  .writedata
		.accelerometer_avalon_accelerometer_spi_mode_slave_byteenable  (mm_interconnect_0_accelerometer_avalon_accelerometer_spi_mode_slave_byteenable),  //                                                  .byteenable
		.accelerometer_avalon_accelerometer_spi_mode_slave_waitrequest (mm_interconnect_0_accelerometer_avalon_accelerometer_spi_mode_slave_waitrequest), //                                                  .waitrequest
		.dram_controller_s1_address                                    (mm_interconnect_0_dram_controller_s1_address),                                    //                                dram_controller_s1.address
		.dram_controller_s1_write                                      (mm_interconnect_0_dram_controller_s1_write),                                      //                                                  .write
		.dram_controller_s1_read                                       (mm_interconnect_0_dram_controller_s1_read),                                       //                                                  .read
		.dram_controller_s1_readdata                                   (mm_interconnect_0_dram_controller_s1_readdata),                                   //                                                  .readdata
		.dram_controller_s1_writedata                                  (mm_interconnect_0_dram_controller_s1_writedata),                                  //                                                  .writedata
		.dram_controller_s1_byteenable                                 (mm_interconnect_0_dram_controller_s1_byteenable),                                 //                                                  .byteenable
		.dram_controller_s1_readdatavalid                              (mm_interconnect_0_dram_controller_s1_readdatavalid),                              //                                                  .readdatavalid
		.dram_controller_s1_waitrequest                                (mm_interconnect_0_dram_controller_s1_waitrequest),                                //                                                  .waitrequest
		.dram_controller_s1_chipselect                                 (mm_interconnect_0_dram_controller_s1_chipselect),                                 //                                                  .chipselect
		.esp32_spi_spi_control_port_address                            (mm_interconnect_0_esp32_spi_spi_control_port_address),                            //                        esp32_spi_spi_control_port.address
		.esp32_spi_spi_control_port_write                              (mm_interconnect_0_esp32_spi_spi_control_port_write),                              //                                                  .write
		.esp32_spi_spi_control_port_read                               (mm_interconnect_0_esp32_spi_spi_control_port_read),                               //                                                  .read
		.esp32_spi_spi_control_port_readdata                           (mm_interconnect_0_esp32_spi_spi_control_port_readdata),                           //                                                  .readdata
		.esp32_spi_spi_control_port_writedata                          (mm_interconnect_0_esp32_spi_spi_control_port_writedata),                          //                                                  .writedata
		.esp32_spi_spi_control_port_chipselect                         (mm_interconnect_0_esp32_spi_spi_control_port_chipselect),                         //                                                  .chipselect
		.jtag_avalon_jtag_slave_address                                (mm_interconnect_0_jtag_avalon_jtag_slave_address),                                //                            jtag_avalon_jtag_slave.address
		.jtag_avalon_jtag_slave_write                                  (mm_interconnect_0_jtag_avalon_jtag_slave_write),                                  //                                                  .write
		.jtag_avalon_jtag_slave_read                                   (mm_interconnect_0_jtag_avalon_jtag_slave_read),                                   //                                                  .read
		.jtag_avalon_jtag_slave_readdata                               (mm_interconnect_0_jtag_avalon_jtag_slave_readdata),                               //                                                  .readdata
		.jtag_avalon_jtag_slave_writedata                              (mm_interconnect_0_jtag_avalon_jtag_slave_writedata),                              //                                                  .writedata
		.jtag_avalon_jtag_slave_waitrequest                            (mm_interconnect_0_jtag_avalon_jtag_slave_waitrequest),                            //                                                  .waitrequest
		.jtag_avalon_jtag_slave_chipselect                             (mm_interconnect_0_jtag_avalon_jtag_slave_chipselect),                             //                                                  .chipselect
		.nios2_cpu_debug_mem_slave_address                             (mm_interconnect_0_nios2_cpu_debug_mem_slave_address),                             //                         nios2_cpu_debug_mem_slave.address
		.nios2_cpu_debug_mem_slave_write                               (mm_interconnect_0_nios2_cpu_debug_mem_slave_write),                               //                                                  .write
		.nios2_cpu_debug_mem_slave_read                                (mm_interconnect_0_nios2_cpu_debug_mem_slave_read),                                //                                                  .read
		.nios2_cpu_debug_mem_slave_readdata                            (mm_interconnect_0_nios2_cpu_debug_mem_slave_readdata),                            //                                                  .readdata
		.nios2_cpu_debug_mem_slave_writedata                           (mm_interconnect_0_nios2_cpu_debug_mem_slave_writedata),                           //                                                  .writedata
		.nios2_cpu_debug_mem_slave_byteenable                          (mm_interconnect_0_nios2_cpu_debug_mem_slave_byteenable),                          //                                                  .byteenable
		.nios2_cpu_debug_mem_slave_waitrequest                         (mm_interconnect_0_nios2_cpu_debug_mem_slave_waitrequest),                         //                                                  .waitrequest
		.nios2_cpu_debug_mem_slave_debugaccess                         (mm_interconnect_0_nios2_cpu_debug_mem_slave_debugaccess),                         //                                                  .debugaccess
		.sys_clk_s1_address                                            (mm_interconnect_0_sys_clk_s1_address),                                            //                                        sys_clk_s1.address
		.sys_clk_s1_write                                              (mm_interconnect_0_sys_clk_s1_write),                                              //                                                  .write
		.sys_clk_s1_readdata                                           (mm_interconnect_0_sys_clk_s1_readdata),                                           //                                                  .readdata
		.sys_clk_s1_writedata                                          (mm_interconnect_0_sys_clk_s1_writedata),                                          //                                                  .writedata
		.sys_clk_s1_chipselect                                         (mm_interconnect_0_sys_clk_s1_chipselect),                                         //                                                  .chipselect
		.timer_1_s1_address                                            (mm_interconnect_0_timer_1_s1_address),                                            //                                        timer_1_s1.address
		.timer_1_s1_write                                              (mm_interconnect_0_timer_1_s1_write),                                              //                                                  .write
		.timer_1_s1_readdata                                           (mm_interconnect_0_timer_1_s1_readdata),                                           //                                                  .readdata
		.timer_1_s1_writedata                                          (mm_interconnect_0_timer_1_s1_writedata),                                          //                                                  .writedata
		.timer_1_s1_chipselect                                         (mm_interconnect_0_timer_1_s1_chipselect),                                         //                                                  .chipselect
		.timer_2_s1_address                                            (mm_interconnect_0_timer_2_s1_address),                                            //                                        timer_2_s1.address
		.timer_2_s1_write                                              (mm_interconnect_0_timer_2_s1_write),                                              //                                                  .write
		.timer_2_s1_readdata                                           (mm_interconnect_0_timer_2_s1_readdata),                                           //                                                  .readdata
		.timer_2_s1_writedata                                          (mm_interconnect_0_timer_2_s1_writedata),                                          //                                                  .writedata
		.timer_2_s1_chipselect                                         (mm_interconnect_0_timer_2_s1_chipselect)                                          //                                                  .chipselect
	);

	esp32SPIHardware_irq_mapper irq_mapper (
		.clk           (dram_clks_pll_sys_clk_clk),      //       clk.clk
		.reset         (rst_controller_reset_out_reset), // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq),       // receiver0.irq
		.receiver1_irq (irq_mapper_receiver1_irq),       // receiver1.irq
		.receiver2_irq (irq_mapper_receiver2_irq),       // receiver2.irq
		.receiver3_irq (irq_mapper_receiver3_irq),       // receiver3.irq
		.receiver4_irq (irq_mapper_receiver4_irq),       // receiver4.irq
		.receiver5_irq (irq_mapper_receiver5_irq),       // receiver5.irq
		.sender_irq    (nios2_cpu_irq_irq)               //    sender.irq
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (dram_clks_pll_reset_source_reset),   // reset_in0.reset
		.clk            (dram_clks_pll_sys_clk_clk),          //       clk.clk
		.reset_out      (rst_controller_reset_out_reset),     // reset_out.reset
		.reset_req      (rst_controller_reset_out_reset_req), //          .reset_req
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_in1      (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_001 (
		.reset_in0      (~reset_reset_n),                     // reset_in0.reset
		.clk            (clk_clk),                            //       clk.clk
		.reset_out      (rst_controller_001_reset_out_reset), // reset_out.reset
		.reset_req      (),                                   // (terminated)
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_in1      (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

endmodule
