// cpu.v

// Generated using ACDS version 20.1 711

`timescale 1 ps / 1 ps
module cpu (
		inout  wire        accelerometer_I2C_SDAT,      // accelerometer.I2C_SDAT
		output wire        accelerometer_I2C_SCLK,      //              .I2C_SCLK
		output wire        accelerometer_G_SENSOR_CS_N, //              .G_SENSOR_CS_N
		input  wire        accelerometer_G_SENSOR_INT,  //              .G_SENSOR_INT
		input  wire        clk_clk,                     //           clk.clk
		output wire [12:0] dram_addr,                   //          dram.addr
		output wire [1:0]  dram_ba,                     //              .ba
		output wire        dram_cas_n,                  //              .cas_n
		output wire        dram_cke,                    //              .cke
		output wire        dram_cs_n,                   //              .cs_n
		inout  wire [15:0] dram_dq,                     //              .dq
		output wire [1:0]  dram_dqm,                    //              .dqm
		output wire        dram_ras_n,                  //              .ras_n
		output wire        dram_we_n,                   //              .we_n
		input  wire        reset_reset_n,               //         reset.reset_n
		output wire        sdram_clk_clk                //     sdram_clk.clk
	);

	wire         pll_sys_clk_clk;                                                                 // pll:sys_clk_clk -> [accelerometer:clk, cpu:clk, integrator_2_0:clk, irq_mapper:clk, jtag:clk, mm_interconnect_0:pll_sys_clk_clk, rst_controller:clk, sdram:clk, timer_0:clk, timer_1:clk]
	wire         cpu_custom_instruction_master_readra;                                            // cpu:D_ci_readra -> cpu_custom_instruction_master_translator:ci_slave_readra
	wire   [4:0] cpu_custom_instruction_master_a;                                                 // cpu:D_ci_a -> cpu_custom_instruction_master_translator:ci_slave_a
	wire   [4:0] cpu_custom_instruction_master_b;                                                 // cpu:D_ci_b -> cpu_custom_instruction_master_translator:ci_slave_b
	wire   [4:0] cpu_custom_instruction_master_c;                                                 // cpu:D_ci_c -> cpu_custom_instruction_master_translator:ci_slave_c
	wire         cpu_custom_instruction_master_readrb;                                            // cpu:D_ci_readrb -> cpu_custom_instruction_master_translator:ci_slave_readrb
	wire         cpu_custom_instruction_master_clk;                                               // cpu:E_ci_multi_clock -> cpu_custom_instruction_master_translator:ci_slave_multi_clk
	wire  [31:0] cpu_custom_instruction_master_ipending;                                          // cpu:W_ci_ipending -> cpu_custom_instruction_master_translator:ci_slave_ipending
	wire         cpu_custom_instruction_master_start;                                             // cpu:E_ci_multi_start -> cpu_custom_instruction_master_translator:ci_slave_multi_start
	wire         cpu_custom_instruction_master_reset_req;                                         // cpu:E_ci_multi_reset_req -> cpu_custom_instruction_master_translator:ci_slave_multi_reset_req
	wire         cpu_custom_instruction_master_done;                                              // cpu_custom_instruction_master_translator:ci_slave_multi_done -> cpu:E_ci_multi_done
	wire   [7:0] cpu_custom_instruction_master_n;                                                 // cpu:D_ci_n -> cpu_custom_instruction_master_translator:ci_slave_n
	wire  [31:0] cpu_custom_instruction_master_result;                                            // cpu_custom_instruction_master_translator:ci_slave_result -> cpu:E_ci_result
	wire         cpu_custom_instruction_master_estatus;                                           // cpu:W_ci_estatus -> cpu_custom_instruction_master_translator:ci_slave_estatus
	wire         cpu_custom_instruction_master_clk_en;                                            // cpu:E_ci_multi_clk_en -> cpu_custom_instruction_master_translator:ci_slave_multi_clken
	wire  [31:0] cpu_custom_instruction_master_datab;                                             // cpu:E_ci_datab -> cpu_custom_instruction_master_translator:ci_slave_datab
	wire  [31:0] cpu_custom_instruction_master_dataa;                                             // cpu:E_ci_dataa -> cpu_custom_instruction_master_translator:ci_slave_dataa
	wire         cpu_custom_instruction_master_reset;                                             // cpu:E_ci_multi_reset -> cpu_custom_instruction_master_translator:ci_slave_multi_reset
	wire         cpu_custom_instruction_master_writerc;                                           // cpu:D_ci_writerc -> cpu_custom_instruction_master_translator:ci_slave_writerc
	wire  [31:0] cpu_custom_instruction_master_translator_comb_ci_master_result;                  // cpu_custom_instruction_master_comb_xconnect:ci_slave_result -> cpu_custom_instruction_master_translator:comb_ci_master_result
	wire         cpu_custom_instruction_master_translator_comb_ci_master_readra;                  // cpu_custom_instruction_master_translator:comb_ci_master_readra -> cpu_custom_instruction_master_comb_xconnect:ci_slave_readra
	wire   [4:0] cpu_custom_instruction_master_translator_comb_ci_master_a;                       // cpu_custom_instruction_master_translator:comb_ci_master_a -> cpu_custom_instruction_master_comb_xconnect:ci_slave_a
	wire   [4:0] cpu_custom_instruction_master_translator_comb_ci_master_b;                       // cpu_custom_instruction_master_translator:comb_ci_master_b -> cpu_custom_instruction_master_comb_xconnect:ci_slave_b
	wire         cpu_custom_instruction_master_translator_comb_ci_master_readrb;                  // cpu_custom_instruction_master_translator:comb_ci_master_readrb -> cpu_custom_instruction_master_comb_xconnect:ci_slave_readrb
	wire   [4:0] cpu_custom_instruction_master_translator_comb_ci_master_c;                       // cpu_custom_instruction_master_translator:comb_ci_master_c -> cpu_custom_instruction_master_comb_xconnect:ci_slave_c
	wire         cpu_custom_instruction_master_translator_comb_ci_master_estatus;                 // cpu_custom_instruction_master_translator:comb_ci_master_estatus -> cpu_custom_instruction_master_comb_xconnect:ci_slave_estatus
	wire  [31:0] cpu_custom_instruction_master_translator_comb_ci_master_ipending;                // cpu_custom_instruction_master_translator:comb_ci_master_ipending -> cpu_custom_instruction_master_comb_xconnect:ci_slave_ipending
	wire  [31:0] cpu_custom_instruction_master_translator_comb_ci_master_datab;                   // cpu_custom_instruction_master_translator:comb_ci_master_datab -> cpu_custom_instruction_master_comb_xconnect:ci_slave_datab
	wire  [31:0] cpu_custom_instruction_master_translator_comb_ci_master_dataa;                   // cpu_custom_instruction_master_translator:comb_ci_master_dataa -> cpu_custom_instruction_master_comb_xconnect:ci_slave_dataa
	wire         cpu_custom_instruction_master_translator_comb_ci_master_writerc;                 // cpu_custom_instruction_master_translator:comb_ci_master_writerc -> cpu_custom_instruction_master_comb_xconnect:ci_slave_writerc
	wire   [7:0] cpu_custom_instruction_master_translator_comb_ci_master_n;                       // cpu_custom_instruction_master_translator:comb_ci_master_n -> cpu_custom_instruction_master_comb_xconnect:ci_slave_n
	wire  [31:0] cpu_custom_instruction_master_comb_xconnect_ci_master0_result;                   // cpu_custom_instruction_master_comb_slave_translator0:ci_slave_result -> cpu_custom_instruction_master_comb_xconnect:ci_master0_result
	wire         cpu_custom_instruction_master_comb_xconnect_ci_master0_readra;                   // cpu_custom_instruction_master_comb_xconnect:ci_master0_readra -> cpu_custom_instruction_master_comb_slave_translator0:ci_slave_readra
	wire   [4:0] cpu_custom_instruction_master_comb_xconnect_ci_master0_a;                        // cpu_custom_instruction_master_comb_xconnect:ci_master0_a -> cpu_custom_instruction_master_comb_slave_translator0:ci_slave_a
	wire   [4:0] cpu_custom_instruction_master_comb_xconnect_ci_master0_b;                        // cpu_custom_instruction_master_comb_xconnect:ci_master0_b -> cpu_custom_instruction_master_comb_slave_translator0:ci_slave_b
	wire         cpu_custom_instruction_master_comb_xconnect_ci_master0_readrb;                   // cpu_custom_instruction_master_comb_xconnect:ci_master0_readrb -> cpu_custom_instruction_master_comb_slave_translator0:ci_slave_readrb
	wire   [4:0] cpu_custom_instruction_master_comb_xconnect_ci_master0_c;                        // cpu_custom_instruction_master_comb_xconnect:ci_master0_c -> cpu_custom_instruction_master_comb_slave_translator0:ci_slave_c
	wire         cpu_custom_instruction_master_comb_xconnect_ci_master0_estatus;                  // cpu_custom_instruction_master_comb_xconnect:ci_master0_estatus -> cpu_custom_instruction_master_comb_slave_translator0:ci_slave_estatus
	wire  [31:0] cpu_custom_instruction_master_comb_xconnect_ci_master0_ipending;                 // cpu_custom_instruction_master_comb_xconnect:ci_master0_ipending -> cpu_custom_instruction_master_comb_slave_translator0:ci_slave_ipending
	wire  [31:0] cpu_custom_instruction_master_comb_xconnect_ci_master0_datab;                    // cpu_custom_instruction_master_comb_xconnect:ci_master0_datab -> cpu_custom_instruction_master_comb_slave_translator0:ci_slave_datab
	wire  [31:0] cpu_custom_instruction_master_comb_xconnect_ci_master0_dataa;                    // cpu_custom_instruction_master_comb_xconnect:ci_master0_dataa -> cpu_custom_instruction_master_comb_slave_translator0:ci_slave_dataa
	wire         cpu_custom_instruction_master_comb_xconnect_ci_master0_writerc;                  // cpu_custom_instruction_master_comb_xconnect:ci_master0_writerc -> cpu_custom_instruction_master_comb_slave_translator0:ci_slave_writerc
	wire   [7:0] cpu_custom_instruction_master_comb_xconnect_ci_master0_n;                        // cpu_custom_instruction_master_comb_xconnect:ci_master0_n -> cpu_custom_instruction_master_comb_slave_translator0:ci_slave_n
	wire  [31:0] cpu_custom_instruction_master_comb_slave_translator0_ci_master_result;           // integrator_2_0:result -> cpu_custom_instruction_master_comb_slave_translator0:ci_master_result
	wire  [31:0] cpu_custom_instruction_master_comb_slave_translator0_ci_master_datab;            // cpu_custom_instruction_master_comb_slave_translator0:ci_master_datab -> integrator_2_0:datab
	wire  [31:0] cpu_custom_instruction_master_comb_slave_translator0_ci_master_dataa;            // cpu_custom_instruction_master_comb_slave_translator0:ci_master_dataa -> integrator_2_0:dataa
	wire  [31:0] cpu_custom_instruction_master_comb_xconnect_ci_master1_result;                   // cpu_custom_instruction_master_comb_slave_translator1:ci_slave_result -> cpu_custom_instruction_master_comb_xconnect:ci_master1_result
	wire         cpu_custom_instruction_master_comb_xconnect_ci_master1_readra;                   // cpu_custom_instruction_master_comb_xconnect:ci_master1_readra -> cpu_custom_instruction_master_comb_slave_translator1:ci_slave_readra
	wire   [4:0] cpu_custom_instruction_master_comb_xconnect_ci_master1_a;                        // cpu_custom_instruction_master_comb_xconnect:ci_master1_a -> cpu_custom_instruction_master_comb_slave_translator1:ci_slave_a
	wire   [4:0] cpu_custom_instruction_master_comb_xconnect_ci_master1_b;                        // cpu_custom_instruction_master_comb_xconnect:ci_master1_b -> cpu_custom_instruction_master_comb_slave_translator1:ci_slave_b
	wire         cpu_custom_instruction_master_comb_xconnect_ci_master1_readrb;                   // cpu_custom_instruction_master_comb_xconnect:ci_master1_readrb -> cpu_custom_instruction_master_comb_slave_translator1:ci_slave_readrb
	wire   [4:0] cpu_custom_instruction_master_comb_xconnect_ci_master1_c;                        // cpu_custom_instruction_master_comb_xconnect:ci_master1_c -> cpu_custom_instruction_master_comb_slave_translator1:ci_slave_c
	wire         cpu_custom_instruction_master_comb_xconnect_ci_master1_estatus;                  // cpu_custom_instruction_master_comb_xconnect:ci_master1_estatus -> cpu_custom_instruction_master_comb_slave_translator1:ci_slave_estatus
	wire  [31:0] cpu_custom_instruction_master_comb_xconnect_ci_master1_ipending;                 // cpu_custom_instruction_master_comb_xconnect:ci_master1_ipending -> cpu_custom_instruction_master_comb_slave_translator1:ci_slave_ipending
	wire  [31:0] cpu_custom_instruction_master_comb_xconnect_ci_master1_datab;                    // cpu_custom_instruction_master_comb_xconnect:ci_master1_datab -> cpu_custom_instruction_master_comb_slave_translator1:ci_slave_datab
	wire  [31:0] cpu_custom_instruction_master_comb_xconnect_ci_master1_dataa;                    // cpu_custom_instruction_master_comb_xconnect:ci_master1_dataa -> cpu_custom_instruction_master_comb_slave_translator1:ci_slave_dataa
	wire         cpu_custom_instruction_master_comb_xconnect_ci_master1_writerc;                  // cpu_custom_instruction_master_comb_xconnect:ci_master1_writerc -> cpu_custom_instruction_master_comb_slave_translator1:ci_slave_writerc
	wire   [7:0] cpu_custom_instruction_master_comb_xconnect_ci_master1_n;                        // cpu_custom_instruction_master_comb_xconnect:ci_master1_n -> cpu_custom_instruction_master_comb_slave_translator1:ci_slave_n
	wire  [31:0] cpu_custom_instruction_master_comb_slave_translator1_ci_master_result;           // nios_custom_instr_floating_point_2_0:s1_result -> cpu_custom_instruction_master_comb_slave_translator1:ci_master_result
	wire  [31:0] cpu_custom_instruction_master_comb_slave_translator1_ci_master_datab;            // cpu_custom_instruction_master_comb_slave_translator1:ci_master_datab -> nios_custom_instr_floating_point_2_0:s1_datab
	wire  [31:0] cpu_custom_instruction_master_comb_slave_translator1_ci_master_dataa;            // cpu_custom_instruction_master_comb_slave_translator1:ci_master_dataa -> nios_custom_instr_floating_point_2_0:s1_dataa
	wire   [3:0] cpu_custom_instruction_master_comb_slave_translator1_ci_master_n;                // cpu_custom_instruction_master_comb_slave_translator1:ci_master_n -> nios_custom_instr_floating_point_2_0:s1_n
	wire         cpu_custom_instruction_master_translator_multi_ci_master_readra;                 // cpu_custom_instruction_master_translator:multi_ci_master_readra -> cpu_custom_instruction_master_multi_xconnect:ci_slave_readra
	wire   [4:0] cpu_custom_instruction_master_translator_multi_ci_master_a;                      // cpu_custom_instruction_master_translator:multi_ci_master_a -> cpu_custom_instruction_master_multi_xconnect:ci_slave_a
	wire   [4:0] cpu_custom_instruction_master_translator_multi_ci_master_b;                      // cpu_custom_instruction_master_translator:multi_ci_master_b -> cpu_custom_instruction_master_multi_xconnect:ci_slave_b
	wire         cpu_custom_instruction_master_translator_multi_ci_master_clk;                    // cpu_custom_instruction_master_translator:multi_ci_master_clk -> cpu_custom_instruction_master_multi_xconnect:ci_slave_clk
	wire         cpu_custom_instruction_master_translator_multi_ci_master_readrb;                 // cpu_custom_instruction_master_translator:multi_ci_master_readrb -> cpu_custom_instruction_master_multi_xconnect:ci_slave_readrb
	wire   [4:0] cpu_custom_instruction_master_translator_multi_ci_master_c;                      // cpu_custom_instruction_master_translator:multi_ci_master_c -> cpu_custom_instruction_master_multi_xconnect:ci_slave_c
	wire         cpu_custom_instruction_master_translator_multi_ci_master_start;                  // cpu_custom_instruction_master_translator:multi_ci_master_start -> cpu_custom_instruction_master_multi_xconnect:ci_slave_start
	wire         cpu_custom_instruction_master_translator_multi_ci_master_reset_req;              // cpu_custom_instruction_master_translator:multi_ci_master_reset_req -> cpu_custom_instruction_master_multi_xconnect:ci_slave_reset_req
	wire         cpu_custom_instruction_master_translator_multi_ci_master_done;                   // cpu_custom_instruction_master_multi_xconnect:ci_slave_done -> cpu_custom_instruction_master_translator:multi_ci_master_done
	wire   [7:0] cpu_custom_instruction_master_translator_multi_ci_master_n;                      // cpu_custom_instruction_master_translator:multi_ci_master_n -> cpu_custom_instruction_master_multi_xconnect:ci_slave_n
	wire  [31:0] cpu_custom_instruction_master_translator_multi_ci_master_result;                 // cpu_custom_instruction_master_multi_xconnect:ci_slave_result -> cpu_custom_instruction_master_translator:multi_ci_master_result
	wire         cpu_custom_instruction_master_translator_multi_ci_master_clk_en;                 // cpu_custom_instruction_master_translator:multi_ci_master_clken -> cpu_custom_instruction_master_multi_xconnect:ci_slave_clken
	wire  [31:0] cpu_custom_instruction_master_translator_multi_ci_master_datab;                  // cpu_custom_instruction_master_translator:multi_ci_master_datab -> cpu_custom_instruction_master_multi_xconnect:ci_slave_datab
	wire  [31:0] cpu_custom_instruction_master_translator_multi_ci_master_dataa;                  // cpu_custom_instruction_master_translator:multi_ci_master_dataa -> cpu_custom_instruction_master_multi_xconnect:ci_slave_dataa
	wire         cpu_custom_instruction_master_translator_multi_ci_master_reset;                  // cpu_custom_instruction_master_translator:multi_ci_master_reset -> cpu_custom_instruction_master_multi_xconnect:ci_slave_reset
	wire         cpu_custom_instruction_master_translator_multi_ci_master_writerc;                // cpu_custom_instruction_master_translator:multi_ci_master_writerc -> cpu_custom_instruction_master_multi_xconnect:ci_slave_writerc
	wire         cpu_custom_instruction_master_multi_xconnect_ci_master0_readra;                  // cpu_custom_instruction_master_multi_xconnect:ci_master0_readra -> cpu_custom_instruction_master_multi_slave_translator0:ci_slave_readra
	wire   [4:0] cpu_custom_instruction_master_multi_xconnect_ci_master0_a;                       // cpu_custom_instruction_master_multi_xconnect:ci_master0_a -> cpu_custom_instruction_master_multi_slave_translator0:ci_slave_a
	wire   [4:0] cpu_custom_instruction_master_multi_xconnect_ci_master0_b;                       // cpu_custom_instruction_master_multi_xconnect:ci_master0_b -> cpu_custom_instruction_master_multi_slave_translator0:ci_slave_b
	wire         cpu_custom_instruction_master_multi_xconnect_ci_master0_readrb;                  // cpu_custom_instruction_master_multi_xconnect:ci_master0_readrb -> cpu_custom_instruction_master_multi_slave_translator0:ci_slave_readrb
	wire   [4:0] cpu_custom_instruction_master_multi_xconnect_ci_master0_c;                       // cpu_custom_instruction_master_multi_xconnect:ci_master0_c -> cpu_custom_instruction_master_multi_slave_translator0:ci_slave_c
	wire         cpu_custom_instruction_master_multi_xconnect_ci_master0_clk;                     // cpu_custom_instruction_master_multi_xconnect:ci_master0_clk -> cpu_custom_instruction_master_multi_slave_translator0:ci_slave_clk
	wire  [31:0] cpu_custom_instruction_master_multi_xconnect_ci_master0_ipending;                // cpu_custom_instruction_master_multi_xconnect:ci_master0_ipending -> cpu_custom_instruction_master_multi_slave_translator0:ci_slave_ipending
	wire         cpu_custom_instruction_master_multi_xconnect_ci_master0_start;                   // cpu_custom_instruction_master_multi_xconnect:ci_master0_start -> cpu_custom_instruction_master_multi_slave_translator0:ci_slave_start
	wire         cpu_custom_instruction_master_multi_xconnect_ci_master0_reset_req;               // cpu_custom_instruction_master_multi_xconnect:ci_master0_reset_req -> cpu_custom_instruction_master_multi_slave_translator0:ci_slave_reset_req
	wire         cpu_custom_instruction_master_multi_xconnect_ci_master0_done;                    // cpu_custom_instruction_master_multi_slave_translator0:ci_slave_done -> cpu_custom_instruction_master_multi_xconnect:ci_master0_done
	wire   [7:0] cpu_custom_instruction_master_multi_xconnect_ci_master0_n;                       // cpu_custom_instruction_master_multi_xconnect:ci_master0_n -> cpu_custom_instruction_master_multi_slave_translator0:ci_slave_n
	wire  [31:0] cpu_custom_instruction_master_multi_xconnect_ci_master0_result;                  // cpu_custom_instruction_master_multi_slave_translator0:ci_slave_result -> cpu_custom_instruction_master_multi_xconnect:ci_master0_result
	wire         cpu_custom_instruction_master_multi_xconnect_ci_master0_estatus;                 // cpu_custom_instruction_master_multi_xconnect:ci_master0_estatus -> cpu_custom_instruction_master_multi_slave_translator0:ci_slave_estatus
	wire         cpu_custom_instruction_master_multi_xconnect_ci_master0_clk_en;                  // cpu_custom_instruction_master_multi_xconnect:ci_master0_clken -> cpu_custom_instruction_master_multi_slave_translator0:ci_slave_clken
	wire  [31:0] cpu_custom_instruction_master_multi_xconnect_ci_master0_datab;                   // cpu_custom_instruction_master_multi_xconnect:ci_master0_datab -> cpu_custom_instruction_master_multi_slave_translator0:ci_slave_datab
	wire  [31:0] cpu_custom_instruction_master_multi_xconnect_ci_master0_dataa;                   // cpu_custom_instruction_master_multi_xconnect:ci_master0_dataa -> cpu_custom_instruction_master_multi_slave_translator0:ci_slave_dataa
	wire         cpu_custom_instruction_master_multi_xconnect_ci_master0_reset;                   // cpu_custom_instruction_master_multi_xconnect:ci_master0_reset -> cpu_custom_instruction_master_multi_slave_translator0:ci_slave_reset
	wire         cpu_custom_instruction_master_multi_xconnect_ci_master0_writerc;                 // cpu_custom_instruction_master_multi_xconnect:ci_master0_writerc -> cpu_custom_instruction_master_multi_slave_translator0:ci_slave_writerc
	wire  [31:0] cpu_custom_instruction_master_multi_slave_translator0_ci_master_result;          // nios_custom_instr_floating_point_2_0:s2_result -> cpu_custom_instruction_master_multi_slave_translator0:ci_master_result
	wire         cpu_custom_instruction_master_multi_slave_translator0_ci_master_clk;             // cpu_custom_instruction_master_multi_slave_translator0:ci_master_clk -> nios_custom_instr_floating_point_2_0:s2_clk
	wire         cpu_custom_instruction_master_multi_slave_translator0_ci_master_clk_en;          // cpu_custom_instruction_master_multi_slave_translator0:ci_master_clken -> nios_custom_instr_floating_point_2_0:s2_clk_en
	wire  [31:0] cpu_custom_instruction_master_multi_slave_translator0_ci_master_datab;           // cpu_custom_instruction_master_multi_slave_translator0:ci_master_datab -> nios_custom_instr_floating_point_2_0:s2_datab
	wire  [31:0] cpu_custom_instruction_master_multi_slave_translator0_ci_master_dataa;           // cpu_custom_instruction_master_multi_slave_translator0:ci_master_dataa -> nios_custom_instr_floating_point_2_0:s2_dataa
	wire         cpu_custom_instruction_master_multi_slave_translator0_ci_master_start;           // cpu_custom_instruction_master_multi_slave_translator0:ci_master_start -> nios_custom_instr_floating_point_2_0:s2_start
	wire         cpu_custom_instruction_master_multi_slave_translator0_ci_master_reset;           // cpu_custom_instruction_master_multi_slave_translator0:ci_master_reset -> nios_custom_instr_floating_point_2_0:s2_reset
	wire         cpu_custom_instruction_master_multi_slave_translator0_ci_master_reset_req;       // cpu_custom_instruction_master_multi_slave_translator0:ci_master_reset_req -> nios_custom_instr_floating_point_2_0:s2_reset_req
	wire         cpu_custom_instruction_master_multi_slave_translator0_ci_master_done;            // nios_custom_instr_floating_point_2_0:s2_done -> cpu_custom_instruction_master_multi_slave_translator0:ci_master_done
	wire   [2:0] cpu_custom_instruction_master_multi_slave_translator0_ci_master_n;               // cpu_custom_instruction_master_multi_slave_translator0:ci_master_n -> nios_custom_instr_floating_point_2_0:s2_n
	wire  [31:0] cpu_data_master_readdata;                                                        // mm_interconnect_0:cpu_data_master_readdata -> cpu:d_readdata
	wire         cpu_data_master_waitrequest;                                                     // mm_interconnect_0:cpu_data_master_waitrequest -> cpu:d_waitrequest
	wire         cpu_data_master_debugaccess;                                                     // cpu:debug_mem_slave_debugaccess_to_roms -> mm_interconnect_0:cpu_data_master_debugaccess
	wire  [27:0] cpu_data_master_address;                                                         // cpu:d_address -> mm_interconnect_0:cpu_data_master_address
	wire   [3:0] cpu_data_master_byteenable;                                                      // cpu:d_byteenable -> mm_interconnect_0:cpu_data_master_byteenable
	wire         cpu_data_master_read;                                                            // cpu:d_read -> mm_interconnect_0:cpu_data_master_read
	wire         cpu_data_master_write;                                                           // cpu:d_write -> mm_interconnect_0:cpu_data_master_write
	wire  [31:0] cpu_data_master_writedata;                                                       // cpu:d_writedata -> mm_interconnect_0:cpu_data_master_writedata
	wire  [31:0] cpu_instruction_master_readdata;                                                 // mm_interconnect_0:cpu_instruction_master_readdata -> cpu:i_readdata
	wire         cpu_instruction_master_waitrequest;                                              // mm_interconnect_0:cpu_instruction_master_waitrequest -> cpu:i_waitrequest
	wire  [27:0] cpu_instruction_master_address;                                                  // cpu:i_address -> mm_interconnect_0:cpu_instruction_master_address
	wire         cpu_instruction_master_read;                                                     // cpu:i_read -> mm_interconnect_0:cpu_instruction_master_read
	wire   [7:0] mm_interconnect_0_accelerometer_avalon_accelerometer_spi_mode_slave_readdata;    // accelerometer:readdata -> mm_interconnect_0:accelerometer_avalon_accelerometer_spi_mode_slave_readdata
	wire         mm_interconnect_0_accelerometer_avalon_accelerometer_spi_mode_slave_waitrequest; // accelerometer:waitrequest -> mm_interconnect_0:accelerometer_avalon_accelerometer_spi_mode_slave_waitrequest
	wire   [0:0] mm_interconnect_0_accelerometer_avalon_accelerometer_spi_mode_slave_address;     // mm_interconnect_0:accelerometer_avalon_accelerometer_spi_mode_slave_address -> accelerometer:address
	wire         mm_interconnect_0_accelerometer_avalon_accelerometer_spi_mode_slave_read;        // mm_interconnect_0:accelerometer_avalon_accelerometer_spi_mode_slave_read -> accelerometer:read
	wire   [0:0] mm_interconnect_0_accelerometer_avalon_accelerometer_spi_mode_slave_byteenable;  // mm_interconnect_0:accelerometer_avalon_accelerometer_spi_mode_slave_byteenable -> accelerometer:byteenable
	wire         mm_interconnect_0_accelerometer_avalon_accelerometer_spi_mode_slave_write;       // mm_interconnect_0:accelerometer_avalon_accelerometer_spi_mode_slave_write -> accelerometer:write
	wire   [7:0] mm_interconnect_0_accelerometer_avalon_accelerometer_spi_mode_slave_writedata;   // mm_interconnect_0:accelerometer_avalon_accelerometer_spi_mode_slave_writedata -> accelerometer:writedata
	wire         mm_interconnect_0_jtag_avalon_jtag_slave_chipselect;                             // mm_interconnect_0:jtag_avalon_jtag_slave_chipselect -> jtag:av_chipselect
	wire  [31:0] mm_interconnect_0_jtag_avalon_jtag_slave_readdata;                               // jtag:av_readdata -> mm_interconnect_0:jtag_avalon_jtag_slave_readdata
	wire         mm_interconnect_0_jtag_avalon_jtag_slave_waitrequest;                            // jtag:av_waitrequest -> mm_interconnect_0:jtag_avalon_jtag_slave_waitrequest
	wire   [0:0] mm_interconnect_0_jtag_avalon_jtag_slave_address;                                // mm_interconnect_0:jtag_avalon_jtag_slave_address -> jtag:av_address
	wire         mm_interconnect_0_jtag_avalon_jtag_slave_read;                                   // mm_interconnect_0:jtag_avalon_jtag_slave_read -> jtag:av_read_n
	wire         mm_interconnect_0_jtag_avalon_jtag_slave_write;                                  // mm_interconnect_0:jtag_avalon_jtag_slave_write -> jtag:av_write_n
	wire  [31:0] mm_interconnect_0_jtag_avalon_jtag_slave_writedata;                              // mm_interconnect_0:jtag_avalon_jtag_slave_writedata -> jtag:av_writedata
	wire  [31:0] mm_interconnect_0_cpu_debug_mem_slave_readdata;                                  // cpu:debug_mem_slave_readdata -> mm_interconnect_0:cpu_debug_mem_slave_readdata
	wire         mm_interconnect_0_cpu_debug_mem_slave_waitrequest;                               // cpu:debug_mem_slave_waitrequest -> mm_interconnect_0:cpu_debug_mem_slave_waitrequest
	wire         mm_interconnect_0_cpu_debug_mem_slave_debugaccess;                               // mm_interconnect_0:cpu_debug_mem_slave_debugaccess -> cpu:debug_mem_slave_debugaccess
	wire   [8:0] mm_interconnect_0_cpu_debug_mem_slave_address;                                   // mm_interconnect_0:cpu_debug_mem_slave_address -> cpu:debug_mem_slave_address
	wire         mm_interconnect_0_cpu_debug_mem_slave_read;                                      // mm_interconnect_0:cpu_debug_mem_slave_read -> cpu:debug_mem_slave_read
	wire   [3:0] mm_interconnect_0_cpu_debug_mem_slave_byteenable;                                // mm_interconnect_0:cpu_debug_mem_slave_byteenable -> cpu:debug_mem_slave_byteenable
	wire         mm_interconnect_0_cpu_debug_mem_slave_write;                                     // mm_interconnect_0:cpu_debug_mem_slave_write -> cpu:debug_mem_slave_write
	wire  [31:0] mm_interconnect_0_cpu_debug_mem_slave_writedata;                                 // mm_interconnect_0:cpu_debug_mem_slave_writedata -> cpu:debug_mem_slave_writedata
	wire         mm_interconnect_0_sdram_s1_chipselect;                                           // mm_interconnect_0:sdram_s1_chipselect -> sdram:az_cs
	wire  [15:0] mm_interconnect_0_sdram_s1_readdata;                                             // sdram:za_data -> mm_interconnect_0:sdram_s1_readdata
	wire         mm_interconnect_0_sdram_s1_waitrequest;                                          // sdram:za_waitrequest -> mm_interconnect_0:sdram_s1_waitrequest
	wire  [24:0] mm_interconnect_0_sdram_s1_address;                                              // mm_interconnect_0:sdram_s1_address -> sdram:az_addr
	wire         mm_interconnect_0_sdram_s1_read;                                                 // mm_interconnect_0:sdram_s1_read -> sdram:az_rd_n
	wire   [1:0] mm_interconnect_0_sdram_s1_byteenable;                                           // mm_interconnect_0:sdram_s1_byteenable -> sdram:az_be_n
	wire         mm_interconnect_0_sdram_s1_readdatavalid;                                        // sdram:za_valid -> mm_interconnect_0:sdram_s1_readdatavalid
	wire         mm_interconnect_0_sdram_s1_write;                                                // mm_interconnect_0:sdram_s1_write -> sdram:az_wr_n
	wire  [15:0] mm_interconnect_0_sdram_s1_writedata;                                            // mm_interconnect_0:sdram_s1_writedata -> sdram:az_data
	wire         mm_interconnect_0_timer_0_s1_chipselect;                                         // mm_interconnect_0:timer_0_s1_chipselect -> timer_0:chipselect
	wire  [15:0] mm_interconnect_0_timer_0_s1_readdata;                                           // timer_0:readdata -> mm_interconnect_0:timer_0_s1_readdata
	wire   [2:0] mm_interconnect_0_timer_0_s1_address;                                            // mm_interconnect_0:timer_0_s1_address -> timer_0:address
	wire         mm_interconnect_0_timer_0_s1_write;                                              // mm_interconnect_0:timer_0_s1_write -> timer_0:write_n
	wire  [15:0] mm_interconnect_0_timer_0_s1_writedata;                                          // mm_interconnect_0:timer_0_s1_writedata -> timer_0:writedata
	wire         mm_interconnect_0_timer_1_s1_chipselect;                                         // mm_interconnect_0:timer_1_s1_chipselect -> timer_1:chipselect
	wire  [15:0] mm_interconnect_0_timer_1_s1_readdata;                                           // timer_1:readdata -> mm_interconnect_0:timer_1_s1_readdata
	wire   [2:0] mm_interconnect_0_timer_1_s1_address;                                            // mm_interconnect_0:timer_1_s1_address -> timer_1:address
	wire         mm_interconnect_0_timer_1_s1_write;                                              // mm_interconnect_0:timer_1_s1_write -> timer_1:write_n
	wire  [15:0] mm_interconnect_0_timer_1_s1_writedata;                                          // mm_interconnect_0:timer_1_s1_writedata -> timer_1:writedata
	wire         irq_mapper_receiver0_irq;                                                        // accelerometer:irq -> irq_mapper:receiver0_irq
	wire         irq_mapper_receiver1_irq;                                                        // jtag:av_irq -> irq_mapper:receiver1_irq
	wire         irq_mapper_receiver2_irq;                                                        // timer_0:irq -> irq_mapper:receiver2_irq
	wire         irq_mapper_receiver3_irq;                                                        // timer_1:irq -> irq_mapper:receiver3_irq
	wire  [31:0] cpu_irq_irq;                                                                     // irq_mapper:sender_irq -> cpu:irq
	wire         rst_controller_reset_out_reset;                                                  // rst_controller:reset_out -> [accelerometer:reset, cpu:reset_n, integrator_2_0:reset, irq_mapper:reset, jtag:rst_n, mm_interconnect_0:cpu_reset_reset_bridge_in_reset_reset, rst_translator:in_reset, sdram:reset_n, timer_0:reset_n, timer_1:reset_n]
	wire         rst_controller_reset_out_reset_req;                                              // rst_controller:reset_req -> [cpu:reset_req, rst_translator:reset_req_in]
	wire         rst_controller_001_reset_out_reset;                                              // rst_controller_001:reset_out -> pll:ref_reset_reset

	cpu_accelerometer accelerometer (
		.clk           (pll_sys_clk_clk),                                                                 //                                 clk.clk
		.reset         (rst_controller_reset_out_reset),                                                  //                               reset.reset
		.address       (mm_interconnect_0_accelerometer_avalon_accelerometer_spi_mode_slave_address),     // avalon_accelerometer_spi_mode_slave.address
		.byteenable    (mm_interconnect_0_accelerometer_avalon_accelerometer_spi_mode_slave_byteenable),  //                                    .byteenable
		.read          (mm_interconnect_0_accelerometer_avalon_accelerometer_spi_mode_slave_read),        //                                    .read
		.write         (mm_interconnect_0_accelerometer_avalon_accelerometer_spi_mode_slave_write),       //                                    .write
		.writedata     (mm_interconnect_0_accelerometer_avalon_accelerometer_spi_mode_slave_writedata),   //                                    .writedata
		.readdata      (mm_interconnect_0_accelerometer_avalon_accelerometer_spi_mode_slave_readdata),    //                                    .readdata
		.waitrequest   (mm_interconnect_0_accelerometer_avalon_accelerometer_spi_mode_slave_waitrequest), //                                    .waitrequest
		.irq           (irq_mapper_receiver0_irq),                                                        //                           interrupt.irq
		.I2C_SDAT      (accelerometer_I2C_SDAT),                                                          //                  external_interface.export
		.I2C_SCLK      (accelerometer_I2C_SCLK),                                                          //                                    .export
		.G_SENSOR_CS_N (accelerometer_G_SENSOR_CS_N),                                                     //                                    .export
		.G_SENSOR_INT  (accelerometer_G_SENSOR_INT)                                                       //                                    .export
	);

	cpu_cpu cpu (
		.clk                                 (pll_sys_clk_clk),                                   //                       clk.clk
		.reset_n                             (~rst_controller_reset_out_reset),                   //                     reset.reset_n
		.reset_req                           (rst_controller_reset_out_reset_req),                //                          .reset_req
		.d_address                           (cpu_data_master_address),                           //               data_master.address
		.d_byteenable                        (cpu_data_master_byteenable),                        //                          .byteenable
		.d_read                              (cpu_data_master_read),                              //                          .read
		.d_readdata                          (cpu_data_master_readdata),                          //                          .readdata
		.d_waitrequest                       (cpu_data_master_waitrequest),                       //                          .waitrequest
		.d_write                             (cpu_data_master_write),                             //                          .write
		.d_writedata                         (cpu_data_master_writedata),                         //                          .writedata
		.debug_mem_slave_debugaccess_to_roms (cpu_data_master_debugaccess),                       //                          .debugaccess
		.i_address                           (cpu_instruction_master_address),                    //        instruction_master.address
		.i_read                              (cpu_instruction_master_read),                       //                          .read
		.i_readdata                          (cpu_instruction_master_readdata),                   //                          .readdata
		.i_waitrequest                       (cpu_instruction_master_waitrequest),                //                          .waitrequest
		.irq                                 (cpu_irq_irq),                                       //                       irq.irq
		.debug_reset_request                 (),                                                  //       debug_reset_request.reset
		.debug_mem_slave_address             (mm_interconnect_0_cpu_debug_mem_slave_address),     //           debug_mem_slave.address
		.debug_mem_slave_byteenable          (mm_interconnect_0_cpu_debug_mem_slave_byteenable),  //                          .byteenable
		.debug_mem_slave_debugaccess         (mm_interconnect_0_cpu_debug_mem_slave_debugaccess), //                          .debugaccess
		.debug_mem_slave_read                (mm_interconnect_0_cpu_debug_mem_slave_read),        //                          .read
		.debug_mem_slave_readdata            (mm_interconnect_0_cpu_debug_mem_slave_readdata),    //                          .readdata
		.debug_mem_slave_waitrequest         (mm_interconnect_0_cpu_debug_mem_slave_waitrequest), //                          .waitrequest
		.debug_mem_slave_write               (mm_interconnect_0_cpu_debug_mem_slave_write),       //                          .write
		.debug_mem_slave_writedata           (mm_interconnect_0_cpu_debug_mem_slave_writedata),   //                          .writedata
		.E_ci_multi_done                     (cpu_custom_instruction_master_done),                // custom_instruction_master.done
		.E_ci_multi_clk_en                   (cpu_custom_instruction_master_clk_en),              //                          .clk_en
		.E_ci_multi_start                    (cpu_custom_instruction_master_start),               //                          .start
		.E_ci_result                         (cpu_custom_instruction_master_result),              //                          .result
		.D_ci_a                              (cpu_custom_instruction_master_a),                   //                          .a
		.D_ci_b                              (cpu_custom_instruction_master_b),                   //                          .b
		.D_ci_c                              (cpu_custom_instruction_master_c),                   //                          .c
		.D_ci_n                              (cpu_custom_instruction_master_n),                   //                          .n
		.D_ci_readra                         (cpu_custom_instruction_master_readra),              //                          .readra
		.D_ci_readrb                         (cpu_custom_instruction_master_readrb),              //                          .readrb
		.D_ci_writerc                        (cpu_custom_instruction_master_writerc),             //                          .writerc
		.E_ci_dataa                          (cpu_custom_instruction_master_dataa),               //                          .dataa
		.E_ci_datab                          (cpu_custom_instruction_master_datab),               //                          .datab
		.E_ci_multi_clock                    (cpu_custom_instruction_master_clk),                 //                          .clk
		.E_ci_multi_reset                    (cpu_custom_instruction_master_reset),               //                          .reset
		.E_ci_multi_reset_req                (cpu_custom_instruction_master_reset_req),           //                          .reset_req
		.W_ci_estatus                        (cpu_custom_instruction_master_estatus),             //                          .estatus
		.W_ci_ipending                       (cpu_custom_instruction_master_ipending)             //                          .ipending
	);

	integrator integrator_2_0 (
		.clk    (pll_sys_clk_clk),                                                       //                         clock.clk
		.reset  (rst_controller_reset_out_reset),                                        //                         reset.reset
		.clk_en (),                                                                      // nios_custom_instruction_slave.clk_en
		.start  (),                                                                      //                              .start
		.done   (),                                                                      //                              .done
		.dataa  (cpu_custom_instruction_master_comb_slave_translator0_ci_master_dataa),  //                              .dataa
		.datab  (cpu_custom_instruction_master_comb_slave_translator0_ci_master_datab),  //                              .datab
		.result (cpu_custom_instruction_master_comb_slave_translator0_ci_master_result)  //                              .result
	);

	cpu_jtag jtag (
		.clk            (pll_sys_clk_clk),                                      //               clk.clk
		.rst_n          (~rst_controller_reset_out_reset),                      //             reset.reset_n
		.av_chipselect  (mm_interconnect_0_jtag_avalon_jtag_slave_chipselect),  // avalon_jtag_slave.chipselect
		.av_address     (mm_interconnect_0_jtag_avalon_jtag_slave_address),     //                  .address
		.av_read_n      (~mm_interconnect_0_jtag_avalon_jtag_slave_read),       //                  .read_n
		.av_readdata    (mm_interconnect_0_jtag_avalon_jtag_slave_readdata),    //                  .readdata
		.av_write_n     (~mm_interconnect_0_jtag_avalon_jtag_slave_write),      //                  .write_n
		.av_writedata   (mm_interconnect_0_jtag_avalon_jtag_slave_writedata),   //                  .writedata
		.av_waitrequest (mm_interconnect_0_jtag_avalon_jtag_slave_waitrequest), //                  .waitrequest
		.av_irq         (irq_mapper_receiver1_irq)                              //               irq.irq
	);

	cpu_nios_custom_instr_floating_point_2_0 #(
		.arithmetic_present (1),
		.root_present       (0),
		.conversion_present (1),
		.comparison_present (1)
	) nios_custom_instr_floating_point_2_0 (
		.s1_dataa     (cpu_custom_instruction_master_comb_slave_translator1_ci_master_dataa),      // s1.dataa
		.s1_datab     (cpu_custom_instruction_master_comb_slave_translator1_ci_master_datab),      //   .datab
		.s1_n         (cpu_custom_instruction_master_comb_slave_translator1_ci_master_n),          //   .n
		.s1_result    (cpu_custom_instruction_master_comb_slave_translator1_ci_master_result),     //   .result
		.s2_clk       (cpu_custom_instruction_master_multi_slave_translator0_ci_master_clk),       // s2.clk
		.s2_clk_en    (cpu_custom_instruction_master_multi_slave_translator0_ci_master_clk_en),    //   .clk_en
		.s2_dataa     (cpu_custom_instruction_master_multi_slave_translator0_ci_master_dataa),     //   .dataa
		.s2_datab     (cpu_custom_instruction_master_multi_slave_translator0_ci_master_datab),     //   .datab
		.s2_n         (cpu_custom_instruction_master_multi_slave_translator0_ci_master_n),         //   .n
		.s2_reset     (cpu_custom_instruction_master_multi_slave_translator0_ci_master_reset),     //   .reset
		.s2_reset_req (cpu_custom_instruction_master_multi_slave_translator0_ci_master_reset_req), //   .reset_req
		.s2_start     (cpu_custom_instruction_master_multi_slave_translator0_ci_master_start),     //   .start
		.s2_done      (cpu_custom_instruction_master_multi_slave_translator0_ci_master_done),      //   .done
		.s2_result    (cpu_custom_instruction_master_multi_slave_translator0_ci_master_result)     //   .result
	);

	cpu_pll pll (
		.ref_clk_clk        (clk_clk),                            //      ref_clk.clk
		.ref_reset_reset    (rst_controller_001_reset_out_reset), //    ref_reset.reset
		.sys_clk_clk        (pll_sys_clk_clk),                    //      sys_clk.clk
		.sdram_clk_clk      (sdram_clk_clk),                      //    sdram_clk.clk
		.reset_source_reset ()                                    // reset_source.reset
	);

	cpu_sdram sdram (
		.clk            (pll_sys_clk_clk),                          //   clk.clk
		.reset_n        (~rst_controller_reset_out_reset),          // reset.reset_n
		.az_addr        (mm_interconnect_0_sdram_s1_address),       //    s1.address
		.az_be_n        (~mm_interconnect_0_sdram_s1_byteenable),   //      .byteenable_n
		.az_cs          (mm_interconnect_0_sdram_s1_chipselect),    //      .chipselect
		.az_data        (mm_interconnect_0_sdram_s1_writedata),     //      .writedata
		.az_rd_n        (~mm_interconnect_0_sdram_s1_read),         //      .read_n
		.az_wr_n        (~mm_interconnect_0_sdram_s1_write),        //      .write_n
		.za_data        (mm_interconnect_0_sdram_s1_readdata),      //      .readdata
		.za_valid       (mm_interconnect_0_sdram_s1_readdatavalid), //      .readdatavalid
		.za_waitrequest (mm_interconnect_0_sdram_s1_waitrequest),   //      .waitrequest
		.zs_addr        (dram_addr),                                //  wire.export
		.zs_ba          (dram_ba),                                  //      .export
		.zs_cas_n       (dram_cas_n),                               //      .export
		.zs_cke         (dram_cke),                                 //      .export
		.zs_cs_n        (dram_cs_n),                                //      .export
		.zs_dq          (dram_dq),                                  //      .export
		.zs_dqm         (dram_dqm),                                 //      .export
		.zs_ras_n       (dram_ras_n),                               //      .export
		.zs_we_n        (dram_we_n)                                 //      .export
	);

	cpu_timer_0 timer_0 (
		.clk        (pll_sys_clk_clk),                         //   clk.clk
		.reset_n    (~rst_controller_reset_out_reset),         // reset.reset_n
		.address    (mm_interconnect_0_timer_0_s1_address),    //    s1.address
		.writedata  (mm_interconnect_0_timer_0_s1_writedata),  //      .writedata
		.readdata   (mm_interconnect_0_timer_0_s1_readdata),   //      .readdata
		.chipselect (mm_interconnect_0_timer_0_s1_chipselect), //      .chipselect
		.write_n    (~mm_interconnect_0_timer_0_s1_write),     //      .write_n
		.irq        (irq_mapper_receiver2_irq)                 //   irq.irq
	);

	cpu_timer_0 timer_1 (
		.clk        (pll_sys_clk_clk),                         //   clk.clk
		.reset_n    (~rst_controller_reset_out_reset),         // reset.reset_n
		.address    (mm_interconnect_0_timer_1_s1_address),    //    s1.address
		.writedata  (mm_interconnect_0_timer_1_s1_writedata),  //      .writedata
		.readdata   (mm_interconnect_0_timer_1_s1_readdata),   //      .readdata
		.chipselect (mm_interconnect_0_timer_1_s1_chipselect), //      .chipselect
		.write_n    (~mm_interconnect_0_timer_1_s1_write),     //      .write_n
		.irq        (irq_mapper_receiver3_irq)                 //   irq.irq
	);

	altera_customins_master_translator #(
		.SHARED_COMB_AND_MULTI (1)
	) cpu_custom_instruction_master_translator (
		.ci_slave_dataa            (cpu_custom_instruction_master_dataa),                                //        ci_slave.dataa
		.ci_slave_datab            (cpu_custom_instruction_master_datab),                                //                .datab
		.ci_slave_result           (cpu_custom_instruction_master_result),                               //                .result
		.ci_slave_n                (cpu_custom_instruction_master_n),                                    //                .n
		.ci_slave_readra           (cpu_custom_instruction_master_readra),                               //                .readra
		.ci_slave_readrb           (cpu_custom_instruction_master_readrb),                               //                .readrb
		.ci_slave_writerc          (cpu_custom_instruction_master_writerc),                              //                .writerc
		.ci_slave_a                (cpu_custom_instruction_master_a),                                    //                .a
		.ci_slave_b                (cpu_custom_instruction_master_b),                                    //                .b
		.ci_slave_c                (cpu_custom_instruction_master_c),                                    //                .c
		.ci_slave_ipending         (cpu_custom_instruction_master_ipending),                             //                .ipending
		.ci_slave_estatus          (cpu_custom_instruction_master_estatus),                              //                .estatus
		.ci_slave_multi_clk        (cpu_custom_instruction_master_clk),                                  //                .clk
		.ci_slave_multi_reset      (cpu_custom_instruction_master_reset),                                //                .reset
		.ci_slave_multi_clken      (cpu_custom_instruction_master_clk_en),                               //                .clk_en
		.ci_slave_multi_reset_req  (cpu_custom_instruction_master_reset_req),                            //                .reset_req
		.ci_slave_multi_start      (cpu_custom_instruction_master_start),                                //                .start
		.ci_slave_multi_done       (cpu_custom_instruction_master_done),                                 //                .done
		.comb_ci_master_dataa      (cpu_custom_instruction_master_translator_comb_ci_master_dataa),      //  comb_ci_master.dataa
		.comb_ci_master_datab      (cpu_custom_instruction_master_translator_comb_ci_master_datab),      //                .datab
		.comb_ci_master_result     (cpu_custom_instruction_master_translator_comb_ci_master_result),     //                .result
		.comb_ci_master_n          (cpu_custom_instruction_master_translator_comb_ci_master_n),          //                .n
		.comb_ci_master_readra     (cpu_custom_instruction_master_translator_comb_ci_master_readra),     //                .readra
		.comb_ci_master_readrb     (cpu_custom_instruction_master_translator_comb_ci_master_readrb),     //                .readrb
		.comb_ci_master_writerc    (cpu_custom_instruction_master_translator_comb_ci_master_writerc),    //                .writerc
		.comb_ci_master_a          (cpu_custom_instruction_master_translator_comb_ci_master_a),          //                .a
		.comb_ci_master_b          (cpu_custom_instruction_master_translator_comb_ci_master_b),          //                .b
		.comb_ci_master_c          (cpu_custom_instruction_master_translator_comb_ci_master_c),          //                .c
		.comb_ci_master_ipending   (cpu_custom_instruction_master_translator_comb_ci_master_ipending),   //                .ipending
		.comb_ci_master_estatus    (cpu_custom_instruction_master_translator_comb_ci_master_estatus),    //                .estatus
		.multi_ci_master_clk       (cpu_custom_instruction_master_translator_multi_ci_master_clk),       // multi_ci_master.clk
		.multi_ci_master_reset     (cpu_custom_instruction_master_translator_multi_ci_master_reset),     //                .reset
		.multi_ci_master_clken     (cpu_custom_instruction_master_translator_multi_ci_master_clk_en),    //                .clk_en
		.multi_ci_master_reset_req (cpu_custom_instruction_master_translator_multi_ci_master_reset_req), //                .reset_req
		.multi_ci_master_start     (cpu_custom_instruction_master_translator_multi_ci_master_start),     //                .start
		.multi_ci_master_done      (cpu_custom_instruction_master_translator_multi_ci_master_done),      //                .done
		.multi_ci_master_dataa     (cpu_custom_instruction_master_translator_multi_ci_master_dataa),     //                .dataa
		.multi_ci_master_datab     (cpu_custom_instruction_master_translator_multi_ci_master_datab),     //                .datab
		.multi_ci_master_result    (cpu_custom_instruction_master_translator_multi_ci_master_result),    //                .result
		.multi_ci_master_n         (cpu_custom_instruction_master_translator_multi_ci_master_n),         //                .n
		.multi_ci_master_readra    (cpu_custom_instruction_master_translator_multi_ci_master_readra),    //                .readra
		.multi_ci_master_readrb    (cpu_custom_instruction_master_translator_multi_ci_master_readrb),    //                .readrb
		.multi_ci_master_writerc   (cpu_custom_instruction_master_translator_multi_ci_master_writerc),   //                .writerc
		.multi_ci_master_a         (cpu_custom_instruction_master_translator_multi_ci_master_a),         //                .a
		.multi_ci_master_b         (cpu_custom_instruction_master_translator_multi_ci_master_b),         //                .b
		.multi_ci_master_c         (cpu_custom_instruction_master_translator_multi_ci_master_c),         //                .c
		.ci_slave_multi_dataa      (32'b00000000000000000000000000000000),                               //     (terminated)
		.ci_slave_multi_datab      (32'b00000000000000000000000000000000),                               //     (terminated)
		.ci_slave_multi_result     (),                                                                   //     (terminated)
		.ci_slave_multi_n          (8'b00000000),                                                        //     (terminated)
		.ci_slave_multi_readra     (1'b0),                                                               //     (terminated)
		.ci_slave_multi_readrb     (1'b0),                                                               //     (terminated)
		.ci_slave_multi_writerc    (1'b0),                                                               //     (terminated)
		.ci_slave_multi_a          (5'b00000),                                                           //     (terminated)
		.ci_slave_multi_b          (5'b00000),                                                           //     (terminated)
		.ci_slave_multi_c          (5'b00000)                                                            //     (terminated)
	);

	cpu_cpu_custom_instruction_master_comb_xconnect cpu_custom_instruction_master_comb_xconnect (
		.ci_slave_dataa      (cpu_custom_instruction_master_translator_comb_ci_master_dataa),    //   ci_slave.dataa
		.ci_slave_datab      (cpu_custom_instruction_master_translator_comb_ci_master_datab),    //           .datab
		.ci_slave_result     (cpu_custom_instruction_master_translator_comb_ci_master_result),   //           .result
		.ci_slave_n          (cpu_custom_instruction_master_translator_comb_ci_master_n),        //           .n
		.ci_slave_readra     (cpu_custom_instruction_master_translator_comb_ci_master_readra),   //           .readra
		.ci_slave_readrb     (cpu_custom_instruction_master_translator_comb_ci_master_readrb),   //           .readrb
		.ci_slave_writerc    (cpu_custom_instruction_master_translator_comb_ci_master_writerc),  //           .writerc
		.ci_slave_a          (cpu_custom_instruction_master_translator_comb_ci_master_a),        //           .a
		.ci_slave_b          (cpu_custom_instruction_master_translator_comb_ci_master_b),        //           .b
		.ci_slave_c          (cpu_custom_instruction_master_translator_comb_ci_master_c),        //           .c
		.ci_slave_ipending   (cpu_custom_instruction_master_translator_comb_ci_master_ipending), //           .ipending
		.ci_slave_estatus    (cpu_custom_instruction_master_translator_comb_ci_master_estatus),  //           .estatus
		.ci_master0_dataa    (cpu_custom_instruction_master_comb_xconnect_ci_master0_dataa),     // ci_master0.dataa
		.ci_master0_datab    (cpu_custom_instruction_master_comb_xconnect_ci_master0_datab),     //           .datab
		.ci_master0_result   (cpu_custom_instruction_master_comb_xconnect_ci_master0_result),    //           .result
		.ci_master0_n        (cpu_custom_instruction_master_comb_xconnect_ci_master0_n),         //           .n
		.ci_master0_readra   (cpu_custom_instruction_master_comb_xconnect_ci_master0_readra),    //           .readra
		.ci_master0_readrb   (cpu_custom_instruction_master_comb_xconnect_ci_master0_readrb),    //           .readrb
		.ci_master0_writerc  (cpu_custom_instruction_master_comb_xconnect_ci_master0_writerc),   //           .writerc
		.ci_master0_a        (cpu_custom_instruction_master_comb_xconnect_ci_master0_a),         //           .a
		.ci_master0_b        (cpu_custom_instruction_master_comb_xconnect_ci_master0_b),         //           .b
		.ci_master0_c        (cpu_custom_instruction_master_comb_xconnect_ci_master0_c),         //           .c
		.ci_master0_ipending (cpu_custom_instruction_master_comb_xconnect_ci_master0_ipending),  //           .ipending
		.ci_master0_estatus  (cpu_custom_instruction_master_comb_xconnect_ci_master0_estatus),   //           .estatus
		.ci_master1_dataa    (cpu_custom_instruction_master_comb_xconnect_ci_master1_dataa),     // ci_master1.dataa
		.ci_master1_datab    (cpu_custom_instruction_master_comb_xconnect_ci_master1_datab),     //           .datab
		.ci_master1_result   (cpu_custom_instruction_master_comb_xconnect_ci_master1_result),    //           .result
		.ci_master1_n        (cpu_custom_instruction_master_comb_xconnect_ci_master1_n),         //           .n
		.ci_master1_readra   (cpu_custom_instruction_master_comb_xconnect_ci_master1_readra),    //           .readra
		.ci_master1_readrb   (cpu_custom_instruction_master_comb_xconnect_ci_master1_readrb),    //           .readrb
		.ci_master1_writerc  (cpu_custom_instruction_master_comb_xconnect_ci_master1_writerc),   //           .writerc
		.ci_master1_a        (cpu_custom_instruction_master_comb_xconnect_ci_master1_a),         //           .a
		.ci_master1_b        (cpu_custom_instruction_master_comb_xconnect_ci_master1_b),         //           .b
		.ci_master1_c        (cpu_custom_instruction_master_comb_xconnect_ci_master1_c),         //           .c
		.ci_master1_ipending (cpu_custom_instruction_master_comb_xconnect_ci_master1_ipending),  //           .ipending
		.ci_master1_estatus  (cpu_custom_instruction_master_comb_xconnect_ci_master1_estatus)    //           .estatus
	);

	altera_customins_slave_translator #(
		.N_WIDTH          (8),
		.USE_DONE         (1),
		.NUM_FIXED_CYCLES (0)
	) cpu_custom_instruction_master_comb_slave_translator0 (
		.ci_slave_dataa      (cpu_custom_instruction_master_comb_xconnect_ci_master0_dataa),          //  ci_slave.dataa
		.ci_slave_datab      (cpu_custom_instruction_master_comb_xconnect_ci_master0_datab),          //          .datab
		.ci_slave_result     (cpu_custom_instruction_master_comb_xconnect_ci_master0_result),         //          .result
		.ci_slave_n          (cpu_custom_instruction_master_comb_xconnect_ci_master0_n),              //          .n
		.ci_slave_readra     (cpu_custom_instruction_master_comb_xconnect_ci_master0_readra),         //          .readra
		.ci_slave_readrb     (cpu_custom_instruction_master_comb_xconnect_ci_master0_readrb),         //          .readrb
		.ci_slave_writerc    (cpu_custom_instruction_master_comb_xconnect_ci_master0_writerc),        //          .writerc
		.ci_slave_a          (cpu_custom_instruction_master_comb_xconnect_ci_master0_a),              //          .a
		.ci_slave_b          (cpu_custom_instruction_master_comb_xconnect_ci_master0_b),              //          .b
		.ci_slave_c          (cpu_custom_instruction_master_comb_xconnect_ci_master0_c),              //          .c
		.ci_slave_ipending   (cpu_custom_instruction_master_comb_xconnect_ci_master0_ipending),       //          .ipending
		.ci_slave_estatus    (cpu_custom_instruction_master_comb_xconnect_ci_master0_estatus),        //          .estatus
		.ci_master_dataa     (cpu_custom_instruction_master_comb_slave_translator0_ci_master_dataa),  // ci_master.dataa
		.ci_master_datab     (cpu_custom_instruction_master_comb_slave_translator0_ci_master_datab),  //          .datab
		.ci_master_result    (cpu_custom_instruction_master_comb_slave_translator0_ci_master_result), //          .result
		.ci_master_n         (),                                                                      // (terminated)
		.ci_master_readra    (),                                                                      // (terminated)
		.ci_master_readrb    (),                                                                      // (terminated)
		.ci_master_writerc   (),                                                                      // (terminated)
		.ci_master_a         (),                                                                      // (terminated)
		.ci_master_b         (),                                                                      // (terminated)
		.ci_master_c         (),                                                                      // (terminated)
		.ci_master_ipending  (),                                                                      // (terminated)
		.ci_master_estatus   (),                                                                      // (terminated)
		.ci_master_clk       (),                                                                      // (terminated)
		.ci_master_clken     (),                                                                      // (terminated)
		.ci_master_reset_req (),                                                                      // (terminated)
		.ci_master_reset     (),                                                                      // (terminated)
		.ci_master_start     (),                                                                      // (terminated)
		.ci_master_done      (1'b0),                                                                  // (terminated)
		.ci_slave_clk        (1'b0),                                                                  // (terminated)
		.ci_slave_clken      (1'b0),                                                                  // (terminated)
		.ci_slave_reset_req  (1'b0),                                                                  // (terminated)
		.ci_slave_reset      (1'b0),                                                                  // (terminated)
		.ci_slave_start      (1'b0),                                                                  // (terminated)
		.ci_slave_done       ()                                                                       // (terminated)
	);

	altera_customins_slave_translator #(
		.N_WIDTH          (4),
		.USE_DONE         (0),
		.NUM_FIXED_CYCLES (0)
	) cpu_custom_instruction_master_comb_slave_translator1 (
		.ci_slave_dataa      (cpu_custom_instruction_master_comb_xconnect_ci_master1_dataa),          //  ci_slave.dataa
		.ci_slave_datab      (cpu_custom_instruction_master_comb_xconnect_ci_master1_datab),          //          .datab
		.ci_slave_result     (cpu_custom_instruction_master_comb_xconnect_ci_master1_result),         //          .result
		.ci_slave_n          (cpu_custom_instruction_master_comb_xconnect_ci_master1_n),              //          .n
		.ci_slave_readra     (cpu_custom_instruction_master_comb_xconnect_ci_master1_readra),         //          .readra
		.ci_slave_readrb     (cpu_custom_instruction_master_comb_xconnect_ci_master1_readrb),         //          .readrb
		.ci_slave_writerc    (cpu_custom_instruction_master_comb_xconnect_ci_master1_writerc),        //          .writerc
		.ci_slave_a          (cpu_custom_instruction_master_comb_xconnect_ci_master1_a),              //          .a
		.ci_slave_b          (cpu_custom_instruction_master_comb_xconnect_ci_master1_b),              //          .b
		.ci_slave_c          (cpu_custom_instruction_master_comb_xconnect_ci_master1_c),              //          .c
		.ci_slave_ipending   (cpu_custom_instruction_master_comb_xconnect_ci_master1_ipending),       //          .ipending
		.ci_slave_estatus    (cpu_custom_instruction_master_comb_xconnect_ci_master1_estatus),        //          .estatus
		.ci_master_dataa     (cpu_custom_instruction_master_comb_slave_translator1_ci_master_dataa),  // ci_master.dataa
		.ci_master_datab     (cpu_custom_instruction_master_comb_slave_translator1_ci_master_datab),  //          .datab
		.ci_master_result    (cpu_custom_instruction_master_comb_slave_translator1_ci_master_result), //          .result
		.ci_master_n         (cpu_custom_instruction_master_comb_slave_translator1_ci_master_n),      //          .n
		.ci_master_readra    (),                                                                      // (terminated)
		.ci_master_readrb    (),                                                                      // (terminated)
		.ci_master_writerc   (),                                                                      // (terminated)
		.ci_master_a         (),                                                                      // (terminated)
		.ci_master_b         (),                                                                      // (terminated)
		.ci_master_c         (),                                                                      // (terminated)
		.ci_master_ipending  (),                                                                      // (terminated)
		.ci_master_estatus   (),                                                                      // (terminated)
		.ci_master_clk       (),                                                                      // (terminated)
		.ci_master_clken     (),                                                                      // (terminated)
		.ci_master_reset_req (),                                                                      // (terminated)
		.ci_master_reset     (),                                                                      // (terminated)
		.ci_master_start     (),                                                                      // (terminated)
		.ci_master_done      (1'b0),                                                                  // (terminated)
		.ci_slave_clk        (1'b0),                                                                  // (terminated)
		.ci_slave_clken      (1'b0),                                                                  // (terminated)
		.ci_slave_reset_req  (1'b0),                                                                  // (terminated)
		.ci_slave_reset      (1'b0),                                                                  // (terminated)
		.ci_slave_start      (1'b0),                                                                  // (terminated)
		.ci_slave_done       ()                                                                       // (terminated)
	);

	cpu_cpu_custom_instruction_master_multi_xconnect cpu_custom_instruction_master_multi_xconnect (
		.ci_slave_dataa       (cpu_custom_instruction_master_translator_multi_ci_master_dataa),     //   ci_slave.dataa
		.ci_slave_datab       (cpu_custom_instruction_master_translator_multi_ci_master_datab),     //           .datab
		.ci_slave_result      (cpu_custom_instruction_master_translator_multi_ci_master_result),    //           .result
		.ci_slave_n           (cpu_custom_instruction_master_translator_multi_ci_master_n),         //           .n
		.ci_slave_readra      (cpu_custom_instruction_master_translator_multi_ci_master_readra),    //           .readra
		.ci_slave_readrb      (cpu_custom_instruction_master_translator_multi_ci_master_readrb),    //           .readrb
		.ci_slave_writerc     (cpu_custom_instruction_master_translator_multi_ci_master_writerc),   //           .writerc
		.ci_slave_a           (cpu_custom_instruction_master_translator_multi_ci_master_a),         //           .a
		.ci_slave_b           (cpu_custom_instruction_master_translator_multi_ci_master_b),         //           .b
		.ci_slave_c           (cpu_custom_instruction_master_translator_multi_ci_master_c),         //           .c
		.ci_slave_ipending    (),                                                                   //           .ipending
		.ci_slave_estatus     (),                                                                   //           .estatus
		.ci_slave_clk         (cpu_custom_instruction_master_translator_multi_ci_master_clk),       //           .clk
		.ci_slave_reset       (cpu_custom_instruction_master_translator_multi_ci_master_reset),     //           .reset
		.ci_slave_clken       (cpu_custom_instruction_master_translator_multi_ci_master_clk_en),    //           .clk_en
		.ci_slave_reset_req   (cpu_custom_instruction_master_translator_multi_ci_master_reset_req), //           .reset_req
		.ci_slave_start       (cpu_custom_instruction_master_translator_multi_ci_master_start),     //           .start
		.ci_slave_done        (cpu_custom_instruction_master_translator_multi_ci_master_done),      //           .done
		.ci_master0_dataa     (cpu_custom_instruction_master_multi_xconnect_ci_master0_dataa),      // ci_master0.dataa
		.ci_master0_datab     (cpu_custom_instruction_master_multi_xconnect_ci_master0_datab),      //           .datab
		.ci_master0_result    (cpu_custom_instruction_master_multi_xconnect_ci_master0_result),     //           .result
		.ci_master0_n         (cpu_custom_instruction_master_multi_xconnect_ci_master0_n),          //           .n
		.ci_master0_readra    (cpu_custom_instruction_master_multi_xconnect_ci_master0_readra),     //           .readra
		.ci_master0_readrb    (cpu_custom_instruction_master_multi_xconnect_ci_master0_readrb),     //           .readrb
		.ci_master0_writerc   (cpu_custom_instruction_master_multi_xconnect_ci_master0_writerc),    //           .writerc
		.ci_master0_a         (cpu_custom_instruction_master_multi_xconnect_ci_master0_a),          //           .a
		.ci_master0_b         (cpu_custom_instruction_master_multi_xconnect_ci_master0_b),          //           .b
		.ci_master0_c         (cpu_custom_instruction_master_multi_xconnect_ci_master0_c),          //           .c
		.ci_master0_ipending  (cpu_custom_instruction_master_multi_xconnect_ci_master0_ipending),   //           .ipending
		.ci_master0_estatus   (cpu_custom_instruction_master_multi_xconnect_ci_master0_estatus),    //           .estatus
		.ci_master0_clk       (cpu_custom_instruction_master_multi_xconnect_ci_master0_clk),        //           .clk
		.ci_master0_reset     (cpu_custom_instruction_master_multi_xconnect_ci_master0_reset),      //           .reset
		.ci_master0_clken     (cpu_custom_instruction_master_multi_xconnect_ci_master0_clk_en),     //           .clk_en
		.ci_master0_reset_req (cpu_custom_instruction_master_multi_xconnect_ci_master0_reset_req),  //           .reset_req
		.ci_master0_start     (cpu_custom_instruction_master_multi_xconnect_ci_master0_start),      //           .start
		.ci_master0_done      (cpu_custom_instruction_master_multi_xconnect_ci_master0_done)        //           .done
	);

	altera_customins_slave_translator #(
		.N_WIDTH          (3),
		.USE_DONE         (1),
		.NUM_FIXED_CYCLES (1)
	) cpu_custom_instruction_master_multi_slave_translator0 (
		.ci_slave_dataa      (cpu_custom_instruction_master_multi_xconnect_ci_master0_dataa),             //  ci_slave.dataa
		.ci_slave_datab      (cpu_custom_instruction_master_multi_xconnect_ci_master0_datab),             //          .datab
		.ci_slave_result     (cpu_custom_instruction_master_multi_xconnect_ci_master0_result),            //          .result
		.ci_slave_n          (cpu_custom_instruction_master_multi_xconnect_ci_master0_n),                 //          .n
		.ci_slave_readra     (cpu_custom_instruction_master_multi_xconnect_ci_master0_readra),            //          .readra
		.ci_slave_readrb     (cpu_custom_instruction_master_multi_xconnect_ci_master0_readrb),            //          .readrb
		.ci_slave_writerc    (cpu_custom_instruction_master_multi_xconnect_ci_master0_writerc),           //          .writerc
		.ci_slave_a          (cpu_custom_instruction_master_multi_xconnect_ci_master0_a),                 //          .a
		.ci_slave_b          (cpu_custom_instruction_master_multi_xconnect_ci_master0_b),                 //          .b
		.ci_slave_c          (cpu_custom_instruction_master_multi_xconnect_ci_master0_c),                 //          .c
		.ci_slave_ipending   (cpu_custom_instruction_master_multi_xconnect_ci_master0_ipending),          //          .ipending
		.ci_slave_estatus    (cpu_custom_instruction_master_multi_xconnect_ci_master0_estatus),           //          .estatus
		.ci_slave_clk        (cpu_custom_instruction_master_multi_xconnect_ci_master0_clk),               //          .clk
		.ci_slave_clken      (cpu_custom_instruction_master_multi_xconnect_ci_master0_clk_en),            //          .clk_en
		.ci_slave_reset_req  (cpu_custom_instruction_master_multi_xconnect_ci_master0_reset_req),         //          .reset_req
		.ci_slave_reset      (cpu_custom_instruction_master_multi_xconnect_ci_master0_reset),             //          .reset
		.ci_slave_start      (cpu_custom_instruction_master_multi_xconnect_ci_master0_start),             //          .start
		.ci_slave_done       (cpu_custom_instruction_master_multi_xconnect_ci_master0_done),              //          .done
		.ci_master_dataa     (cpu_custom_instruction_master_multi_slave_translator0_ci_master_dataa),     // ci_master.dataa
		.ci_master_datab     (cpu_custom_instruction_master_multi_slave_translator0_ci_master_datab),     //          .datab
		.ci_master_result    (cpu_custom_instruction_master_multi_slave_translator0_ci_master_result),    //          .result
		.ci_master_n         (cpu_custom_instruction_master_multi_slave_translator0_ci_master_n),         //          .n
		.ci_master_clk       (cpu_custom_instruction_master_multi_slave_translator0_ci_master_clk),       //          .clk
		.ci_master_clken     (cpu_custom_instruction_master_multi_slave_translator0_ci_master_clk_en),    //          .clk_en
		.ci_master_reset_req (cpu_custom_instruction_master_multi_slave_translator0_ci_master_reset_req), //          .reset_req
		.ci_master_reset     (cpu_custom_instruction_master_multi_slave_translator0_ci_master_reset),     //          .reset
		.ci_master_start     (cpu_custom_instruction_master_multi_slave_translator0_ci_master_start),     //          .start
		.ci_master_done      (cpu_custom_instruction_master_multi_slave_translator0_ci_master_done),      //          .done
		.ci_master_readra    (),                                                                          // (terminated)
		.ci_master_readrb    (),                                                                          // (terminated)
		.ci_master_writerc   (),                                                                          // (terminated)
		.ci_master_a         (),                                                                          // (terminated)
		.ci_master_b         (),                                                                          // (terminated)
		.ci_master_c         (),                                                                          // (terminated)
		.ci_master_ipending  (),                                                                          // (terminated)
		.ci_master_estatus   ()                                                                           // (terminated)
	);

	cpu_mm_interconnect_0 mm_interconnect_0 (
		.pll_sys_clk_clk                                               (pll_sys_clk_clk),                                                                 //                                       pll_sys_clk.clk
		.cpu_reset_reset_bridge_in_reset_reset                         (rst_controller_reset_out_reset),                                                  //                   cpu_reset_reset_bridge_in_reset.reset
		.cpu_data_master_address                                       (cpu_data_master_address),                                                         //                                   cpu_data_master.address
		.cpu_data_master_waitrequest                                   (cpu_data_master_waitrequest),                                                     //                                                  .waitrequest
		.cpu_data_master_byteenable                                    (cpu_data_master_byteenable),                                                      //                                                  .byteenable
		.cpu_data_master_read                                          (cpu_data_master_read),                                                            //                                                  .read
		.cpu_data_master_readdata                                      (cpu_data_master_readdata),                                                        //                                                  .readdata
		.cpu_data_master_write                                         (cpu_data_master_write),                                                           //                                                  .write
		.cpu_data_master_writedata                                     (cpu_data_master_writedata),                                                       //                                                  .writedata
		.cpu_data_master_debugaccess                                   (cpu_data_master_debugaccess),                                                     //                                                  .debugaccess
		.cpu_instruction_master_address                                (cpu_instruction_master_address),                                                  //                            cpu_instruction_master.address
		.cpu_instruction_master_waitrequest                            (cpu_instruction_master_waitrequest),                                              //                                                  .waitrequest
		.cpu_instruction_master_read                                   (cpu_instruction_master_read),                                                     //                                                  .read
		.cpu_instruction_master_readdata                               (cpu_instruction_master_readdata),                                                 //                                                  .readdata
		.accelerometer_avalon_accelerometer_spi_mode_slave_address     (mm_interconnect_0_accelerometer_avalon_accelerometer_spi_mode_slave_address),     // accelerometer_avalon_accelerometer_spi_mode_slave.address
		.accelerometer_avalon_accelerometer_spi_mode_slave_write       (mm_interconnect_0_accelerometer_avalon_accelerometer_spi_mode_slave_write),       //                                                  .write
		.accelerometer_avalon_accelerometer_spi_mode_slave_read        (mm_interconnect_0_accelerometer_avalon_accelerometer_spi_mode_slave_read),        //                                                  .read
		.accelerometer_avalon_accelerometer_spi_mode_slave_readdata    (mm_interconnect_0_accelerometer_avalon_accelerometer_spi_mode_slave_readdata),    //                                                  .readdata
		.accelerometer_avalon_accelerometer_spi_mode_slave_writedata   (mm_interconnect_0_accelerometer_avalon_accelerometer_spi_mode_slave_writedata),   //                                                  .writedata
		.accelerometer_avalon_accelerometer_spi_mode_slave_byteenable  (mm_interconnect_0_accelerometer_avalon_accelerometer_spi_mode_slave_byteenable),  //                                                  .byteenable
		.accelerometer_avalon_accelerometer_spi_mode_slave_waitrequest (mm_interconnect_0_accelerometer_avalon_accelerometer_spi_mode_slave_waitrequest), //                                                  .waitrequest
		.cpu_debug_mem_slave_address                                   (mm_interconnect_0_cpu_debug_mem_slave_address),                                   //                               cpu_debug_mem_slave.address
		.cpu_debug_mem_slave_write                                     (mm_interconnect_0_cpu_debug_mem_slave_write),                                     //                                                  .write
		.cpu_debug_mem_slave_read                                      (mm_interconnect_0_cpu_debug_mem_slave_read),                                      //                                                  .read
		.cpu_debug_mem_slave_readdata                                  (mm_interconnect_0_cpu_debug_mem_slave_readdata),                                  //                                                  .readdata
		.cpu_debug_mem_slave_writedata                                 (mm_interconnect_0_cpu_debug_mem_slave_writedata),                                 //                                                  .writedata
		.cpu_debug_mem_slave_byteenable                                (mm_interconnect_0_cpu_debug_mem_slave_byteenable),                                //                                                  .byteenable
		.cpu_debug_mem_slave_waitrequest                               (mm_interconnect_0_cpu_debug_mem_slave_waitrequest),                               //                                                  .waitrequest
		.cpu_debug_mem_slave_debugaccess                               (mm_interconnect_0_cpu_debug_mem_slave_debugaccess),                               //                                                  .debugaccess
		.jtag_avalon_jtag_slave_address                                (mm_interconnect_0_jtag_avalon_jtag_slave_address),                                //                            jtag_avalon_jtag_slave.address
		.jtag_avalon_jtag_slave_write                                  (mm_interconnect_0_jtag_avalon_jtag_slave_write),                                  //                                                  .write
		.jtag_avalon_jtag_slave_read                                   (mm_interconnect_0_jtag_avalon_jtag_slave_read),                                   //                                                  .read
		.jtag_avalon_jtag_slave_readdata                               (mm_interconnect_0_jtag_avalon_jtag_slave_readdata),                               //                                                  .readdata
		.jtag_avalon_jtag_slave_writedata                              (mm_interconnect_0_jtag_avalon_jtag_slave_writedata),                              //                                                  .writedata
		.jtag_avalon_jtag_slave_waitrequest                            (mm_interconnect_0_jtag_avalon_jtag_slave_waitrequest),                            //                                                  .waitrequest
		.jtag_avalon_jtag_slave_chipselect                             (mm_interconnect_0_jtag_avalon_jtag_slave_chipselect),                             //                                                  .chipselect
		.sdram_s1_address                                              (mm_interconnect_0_sdram_s1_address),                                              //                                          sdram_s1.address
		.sdram_s1_write                                                (mm_interconnect_0_sdram_s1_write),                                                //                                                  .write
		.sdram_s1_read                                                 (mm_interconnect_0_sdram_s1_read),                                                 //                                                  .read
		.sdram_s1_readdata                                             (mm_interconnect_0_sdram_s1_readdata),                                             //                                                  .readdata
		.sdram_s1_writedata                                            (mm_interconnect_0_sdram_s1_writedata),                                            //                                                  .writedata
		.sdram_s1_byteenable                                           (mm_interconnect_0_sdram_s1_byteenable),                                           //                                                  .byteenable
		.sdram_s1_readdatavalid                                        (mm_interconnect_0_sdram_s1_readdatavalid),                                        //                                                  .readdatavalid
		.sdram_s1_waitrequest                                          (mm_interconnect_0_sdram_s1_waitrequest),                                          //                                                  .waitrequest
		.sdram_s1_chipselect                                           (mm_interconnect_0_sdram_s1_chipselect),                                           //                                                  .chipselect
		.timer_0_s1_address                                            (mm_interconnect_0_timer_0_s1_address),                                            //                                        timer_0_s1.address
		.timer_0_s1_write                                              (mm_interconnect_0_timer_0_s1_write),                                              //                                                  .write
		.timer_0_s1_readdata                                           (mm_interconnect_0_timer_0_s1_readdata),                                           //                                                  .readdata
		.timer_0_s1_writedata                                          (mm_interconnect_0_timer_0_s1_writedata),                                          //                                                  .writedata
		.timer_0_s1_chipselect                                         (mm_interconnect_0_timer_0_s1_chipselect),                                         //                                                  .chipselect
		.timer_1_s1_address                                            (mm_interconnect_0_timer_1_s1_address),                                            //                                        timer_1_s1.address
		.timer_1_s1_write                                              (mm_interconnect_0_timer_1_s1_write),                                              //                                                  .write
		.timer_1_s1_readdata                                           (mm_interconnect_0_timer_1_s1_readdata),                                           //                                                  .readdata
		.timer_1_s1_writedata                                          (mm_interconnect_0_timer_1_s1_writedata),                                          //                                                  .writedata
		.timer_1_s1_chipselect                                         (mm_interconnect_0_timer_1_s1_chipselect)                                          //                                                  .chipselect
	);

	cpu_irq_mapper irq_mapper (
		.clk           (pll_sys_clk_clk),                //       clk.clk
		.reset         (rst_controller_reset_out_reset), // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq),       // receiver0.irq
		.receiver1_irq (irq_mapper_receiver1_irq),       // receiver1.irq
		.receiver2_irq (irq_mapper_receiver2_irq),       // receiver2.irq
		.receiver3_irq (irq_mapper_receiver3_irq),       // receiver3.irq
		.sender_irq    (cpu_irq_irq)                     //    sender.irq
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~reset_reset_n),                     // reset_in0.reset
		.clk            (pll_sys_clk_clk),                    //       clk.clk
		.reset_out      (rst_controller_reset_out_reset),     // reset_out.reset
		.reset_req      (rst_controller_reset_out_reset_req), //          .reset_req
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_in1      (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_001 (
		.reset_in0      (~reset_reset_n),                     // reset_in0.reset
		.clk            (clk_clk),                            //       clk.clk
		.reset_out      (rst_controller_001_reset_out_reset), // reset_out.reset
		.reset_req      (),                                   // (terminated)
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_in1      (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

endmodule
